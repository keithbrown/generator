��     &  _H  _Ww %  C o l o r   C h o o s e r�M��". C o l o r   C h o o s e r   O v e r v i e w V i e w s   M e n u ��� ��  ��   ��   ��   ��   ��   ��      �� 	 �� 
 ��  ����     ����  ��    �� ��  ��  ��  ��   �� ����$ S p e c i f y i n g   C o l o r s. Y) �}����5Ni���4a���  O p t i o n s   M e n u C o l o r   B o x2 C o l o r   M e t h o d   P o p - u p   M e n u S a v e d   C o l o r s  C o l o r   V i e w   A r e a C o l o r   W h e e l C o l o r   P l a n e N a m e d   C o l o r s, C o l o r   T o l e r a n c e s   V i e w8 C o l o r   C o m p o n e n t   S l i d e r   B a r s R e f o r m   S l i d e r s* C o n f i r m a t i o n   B u t t o n s C o l o r   M o d e l s, G r a y s c a l e   C o l o r   M o d e l  H L S   C o l o r   M o d e l  R G B   C o l o r   M o d e l  C M Y   C o l o r   M o d e l" C o l o r   T o l e r a n c e s   &'%$ B D e f a u l t   C o l o r   T o l e r a n c e s   D e t a i l s C o l o r W h e e l4C��$C\o�����9Lcz�����*    *   B I m a g e E d i t o r P a l e d D i a l o g v c o l o r c h s r R G B M o d e l   
	  C M Y M o d e l T o l e r a n c e s V i e w S a v e d C o l o r s O v e r v i e w G r a y s c a l e M o d e l C o l o r S l i d e r s V i e w s M e n u P o p U p M e n u R e f o r m S l i d e r s C o l o r B o x C o l o r M o d e l s S p e c i f y C o l o r s H L S M o d e l T o l e r a n c e s v c o l o r c h s r C o l o r V i e w A r e a O p t i o n s M e n u N a m e d C o l o r s C o l o r P l a n e C o n f i r m B u t t o n s* v s t y l e c h s r v c o l o r c h s r" T o l e r a n c e s D e t a i l c o l o r   c h o o s e r (  #!V3?IV\hq{������������)4*+,-./012 S p e c i f y C o l o r s  --
�    ( S a v e d C o l o r s
�    S� C o l o r   C h o o s e r 
 
 U s e   t h e   C o l o r   C h o o s e r   t o   s p e c i f y   c o l o r s   f o r   a n   a p p l i c a t i o n .   Y o u   c a n   s a v e   s p e c i f i e d   c o l o r s ,   a n d   r e v e r t   t o   a   p r e v i o u s   s e l e c t i o n . 
 
 T h e   C o l o r   C h o o s e r   c o n t a i n s   t h e   f o l l o w i n g   c o m p o n e n t s : 
 
 V i e w s   M e n u 
 O p t i o n s   M e n u 
 C o l o r   M e t h o d   P o p   U p   M e n u 
 C o l o r   V i e w   A r e a   ( C o l o r   W h e e l   o r   P l a n e ) 
 C o l o r   S e l e c t i o n   B o x 
 C o l o r   S l i d e r s 
 S a v e d   C o l o r   P a l e t t e 
 C o n f i r m a t i o n   B u t t o n s 
 
 C o l o r B o x

�    n V i e w s M e n u

� 
   � O p t i o n s M e n u
    � P o p U p M e n u
8    � C o l o r V i e w A r e a
X    � C o l o r B o x
�    C o l o r S l i d e r s
�   1 S a v e d C o l o r s
�   ?
    S  B C o n f i r m B u t t o n s� T o   s p e c i f y   c o l o r s ,   d o   a n y   o f   t h e   f o l l o w i n g : 
 
 * 	 S e l e c t   a   c o l o r   m o d e l   f r o m   t h e   C o l o r   M e t h o d   P o p - u p   M e n u . 
 
 * 	 D r a g   t h e   p o i n t e r   i n   t h e   C o l o r   W h e e l   o r   C o l o r   P l a n e .   
 
 * 	 C l i c k   o n   a   C o l o r   C o m p o n e n t   S l i d e r   B a r   o r   d r a g   i t s   i n d i c a t o r   t o   a   n e w   p o s i t i o n .   Y o u   c a n   a l s o   s p e c i f y   v a l u e s   i n   t h e   p e r c e n t a g e   f i e l d s . 
 
 * 	 D o u b l e - c l i c k   o n   a   s a v e d   c o l o r   o n   t h e   S a v e d   C o l o r   P a l e t t e . 
 
 * 	 R e v e r t   t o   a   p r e v i o u s l y   s e l e c t e d   c o l o r   b y   d o u b l e - c l i c k i n g   i n   t h e   t o p   h a l f   o f   t h e   C o l o r   S e l e c t i o n   B o x . 
 
 
 
 

 + +��7865 9 :@;<=> P o p U p M e n u "  
�    M C o l o r W h e e l
    � C o l o r P l a n e
6    � C o l o r S l i d e r s
X    � S a v e d C o l o r s
~   O C o l o r B o x
�   �o V i e w s   M e n u 
 
 U s e   t h e   V i e w s   M e n u   t o   s e l e c t   o n e   o f   t h e   t h r e e   v i e w s   a v a i l a b l e   f o r   t h e   C o l o r   V i e w   A r e a .   T h e   v i e w s   a v a i l a b l e   a r e : 
 
 C o l o r   W h e e l / C o l o r   P l a n e 
 
 N a m e d   C o l o r s 
 
 C o l o r   T o l e r a n c e s 
 
FJGHCDBA E�  C o l o r W h e e l O  
N    } C o l o r P l a n e
y    � N a m e d C o l o r s
�    � T o l e r a n c e s V i e w
�    �MNLKX "�   C C C ��l|III��   / 9    X X W P P	aaV       00 	PWQRSTU R e f o r m S l i d e r s
] #  k C o l o r P l a n e
�   & C o l o r P l a n e
�    N a m e d C o l o r s
�   �
�   dL�	� O p t i o n s   M e n u 
 
 T h e   O p t i o n s   M e n u   c o n t a i n s   t h e   f o l l o w i n g   m e n u   i t e m s : 
 
 R e f o r m   S l i d e r   I m a g e s 
 U s e   t h i s   o p t i o n   t o   s p e c i f y   t h e   a p p e a r a n c e   a n d   b e h a v i o r   o f   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s . 
 
 R e d - G r e e n   P l a n e 
 R e d - B l u e   P l a n e 
 B l u e - G r e e n   P l a n e 
 T h e s e   m e n u   i t e m s   a r e   e n a b l e d   w h e n   t h e   C o l o r   V i e w   A r e a   d e p i c t s   t h e   R G B   C o l o r   P l a n e .   T h e   s e l e c t e d   v a l u e   i n d i c a t e s   w h i c h   c o l o r   p l a n e   i s   d e p i c t e d   i n   t h e   C o l o r   V i e w   A r e a . 
 
 C y a n - M a g e n t a   P l a n e 
 C y a n - Y e l l o w   P l a n e 
 M a g e n t a - Y e l l o w   P l a n e 
 T h e s e   m e n u   i t e m s   a r e   e n a b l e d   w h e n   t h e   C o l o r   V i e w   A r e a   d e p i c t s   t h e   C M Y   C o l o r   P l a n e .   T h e   s e l e c t e d   v a l u e   i n d i c a t e s   w h i c h   c o l o r   p l a n e   i s   d e p i c t e d   i n   t h e   C o l o r   V i e w   A r e a . 
 
 S o r t   b y   N a m e 
 S o r t   b y   H u e 
 T h e s e   m e n u   i t e m s   a r e   e n a b l e d   w h e n   t h e   C o l o r   V i e w   A r e a   d e p i c t s   N a m e d   C o l o r s .   U s e   t h e s e   o p t i o n s   t o   s p e c i f y   t h e   s o r t i n g   o r d e r   o f   t h e   l i s t   o f   N a m e d   C o l o r s . 
 
 
 A d d   S a v e d   C o l o r 
 U s e   t h i s   m e n u   i t e m   t o   a d d   t h e   s p e c i f i e d   c o l o r   t o   t h e   S a v e d   C o l o r s   P a l e t t e . 
 
 
 D e f a u l t   C o l o r   T o l e r a n c e s 
 U s e   t h i s   o p t i o n   t o   s p e c i f y   t h e   d e f a u l t   c o l o r   t o l e r a n c e s   f o r   s e l e c t e d   c o l o r s .   A l l   s e l e c t e d   c o l o r s   w i l l   b e   r e p r e s e n t e d   w i t h   t h e   s e l e c t e d   c o l o r   t o l e r a n c e .   T h e   c h o i c e s   a v a i l a b l e   a r e : 
 
 L a r g e   D i t h e r 
 S m a l l   D i t h e r 
 S o l i d 
 P r e c i s e   L a r g e   D i t h e r 
 P r e c i s e   S m a l l   D i t h e r 
 P r e c i s e   S o l i d 
 
 Y o u   c a n   a l s o   c h a n g e   t h e   d e f a u l t   c o l o r   t o l e r a n c e s   i n   t h e   C o l o r   T o l e r a n c e s   V i e w . 
 
 S a v e d C o l o r s T o l e r a n c e s
   � T o l e r a n c e s V i e w
#   �Z[YX$^0 _`^] a$  	bicdefg C o l o r M o d e l slmkj 
�    K H L S M o d e l
�    � R G B M o d e l
�    � C M Y M o d e l
�    � G r a y s c a l e M o d e l
 	   � C o l o r V i e w A r e a
6    � C o l o r S l i d e r s
^    �  ==KK8 j	++77221e& n(  orp T o l e r a n c e stL 
�    � O p t i o n s M e n u� T h e   C o l o r   B o x 
 
 T h e   C o l o r   B o x   d i s p l a y s   c o l o r   s e l e c t i o n s   i n   t h e   C o l o r   C h o o s e r . 
 
 T h e   b o t t o m   h a l f   o f   t h e   C o l o r   B o x   d i s p l a y s   t h e   c u r r e n t   c o l o r   s e l e c t i o n .   T h e   t o p   h a l f   o f   t h e   C o l o r   B o x   d i s p l a y s   t h e   p r e v i o u s   c o l o r   s e l e c t i o n . 
 
 Y o u   c a n   r e v e r t   f r o m   t h e   c u r r e n t   c o l o r   s e l e c t i o n   t o   t h e   p r e v i o u s   s e l e c t i o n   b y   c l i c k i n g   i n   t h e   t o p   h a l f   o f   t h e   C o l o r   B o x . 
 

�   � C o l o r B o x
"� 	  uvts w0, x|yz C o l o r W h e e l�~} 
"�    � C o l o r P l a n e
#     � N a m e d C o l o r s
#B    � T o l e r a n c e s V i e w
#f    �

		--   = = E E r rYY 1ef& �4  ����� H L S M o d e l���� 
#�    �44i T h e   C o l o r   M e t h o d   P o p - u p   M e n u 
 
 U s e   t h e   C o l o r   M e t h o d   P o p - u p   M e n u   t o   s e l e c t   a   c o l o r   m o d e l   t o   u s e   w h e n   s p e c i f y i n g   a   c o l o r . 
 
 T h e r e   a r e   f o u r   c o l o r   m o d e l s   t o   c h o o s e   f r o m : 
 
 H L S 
 R G B 
 C M Y 
 G r a y s c a l e 
 
 W h e n   a   C o l o r   M o d e l   i s   s e l e c t e d ,   t h e   C o l o r   V i e w   A r e a   a n d   C o l o r   C o m p o n e n t   S l i d e r   B a r s   c h a n g e   t o   r e f l e c t   y o u r   s e l e c t i o n . 
 
 C o l o r B o x
&j 	  # C o l o r S l i d e r s
&�   � T o l e r a n c e s
&�   � T o l e r a n c e s V i e w
&�   !  ee�1% �@  	���������  R G B M o d e l
''   � C M Y M o d e l
'E   � O p t i o n s M e n u
'c   % C o l o r B o x
'� 	  � C o l o r S l i d e r s
'�   � T o l e r a n c e s
'�   �
>�   &"+ S a v e d   C o l o r s 
 
 U s e   t h e   S a v e d   C o l o r s   P a l e t t e   t o   s a v e   f r e q u e n t l y   u s e d   c o l o r s .   Y o u   c a n   s a v e   u p   t o   1 6   c o l o r s   o n   t h e   S a v e d   C o l o r s   P a l e t t e . 
 
 S a v e d   c o l o r s   a r e   a u t o m a t i c a l l y   s a v e d   w i t h   t h e   C o l o r   C h o o s e r   a n d   a r e   a v a i l a b l e   f o r   f u t u r e   e d i t i n g   s e s s i o n s .   T h e   c o l o r   t o l e r a n c e   v a l u e s   f o r   d i t h e r i n g   a r e   s a v e d   w i t h   t h e   s a v e d   c o l o r s . 
 
 
 T o   S a v e   a   C o l o r   o n   t h e   S a v e d   C o l o r   P a l e t t e : 
 
 1 .   S e l e c t   a   c o l o r   i n   t h e   C o l o r   C h o o s e r . 
 
 2 .   P r e s s   t h e   C o n t r o l   k e y   a n d   c l i c k   o n   a   c e l l   i n   t h e   S a v e d   C o l o r   P a l e t t e . 
 
 T h e   c o l o r   i s   s a v e d   i n   t h e   s e l e c t e d   c e l l . 
 
 
 T o   S a v e   a   C o l o r   o n   t h e   S a v e d   C o l o r   P a l e t t e   ( v e r s i o n   2 ) : 
 
 1 .   S e l e c t   a   c o l o r   i n   t h e   C o l o r   C h o o s e r . 
 
 2 .   C l i c k   o n   t h e   S a v e d   C o l o r s   P a l e t t e ,   a n d   u s e   t h e   a r r o w   k e y s   f r o m   t h e   k e y b o a r d   t o   m o v e   t o   a   c e l l   o n   t h e   p a l e t t e . 
 
 3 .   S e l e c t   A d d   S a v e d   C o l o r   f r o m   t h e   O p t i o n s   M e n u   t o   s a v e   t h e   c o l o r . 
 
 T h e   c o l o r   i s   s a v e d   i n   t h e   s e l e c t e d   c e l l . 
 
 
 T o   r e t r i e v e   a   c o l o r   f r o m   t h e   S a v e d   C o l o r s   P a l e t t e : 
 
 1 .   D o u b l e - c l i c k   o n   a   c e l l   i n   t h e   S a v e d   C o l o r s   P a l e t t e . 
 
 T h e   c o l o r   s t o r e d   i n   t h e   c e l l   i s   n o w   t h e   s e l e c t e d   c o l o r ,   a n d   i s   d i s p l a y e d   i n   t h e   C o l o r   B o x . 
 
 
� T h e   C o l o r   V i e w   A r e a 
 
 T h e   C o l o r   V i e w   A r e a   d i s p l a y s   t o o l s   f o r   s e l e c t i n g   a n d   d e f i n i n g   c o l o r s   f o r   y o u r   a p p l i c a t i o n .   T h r e e   d i f f e r e n t   v i e w s   a r e   a v a i l a b l e : 
 
 C o l o r   W h e e l / C o l o r   P l a n e 
 N a m e d   C o l o r s 
 C o l o r   T o l e r a n c e s 
 
 T h e   C o l o r   W h e e l / C o l o r   P l a n e   v i e w   d i s p l a y s   a   g r a p h i c   r e p r e s e n t a t i o n ,   o r   m a p ,   o f   t h e   s e l e c t e d   c o l o r   m o d e l .   T h e   N a m e d   C o l o r s   v i e w   d i s p l a y s   a   s c r o l l i n g   l i s t   o f   p r e d e f i n e d   c o l o r s .   T h e   C o l o r   T o l e r a n c e s   d i s p l a y s   a   s e t   o f   t o o l s   y o u   c a n   u s e   t o   d e f i n e   t h e   a p p e a r a n c e   o f   c o l o r s   o n   a   d i s p l a y . 
 
 

� T h e   H L S   C o l o r   W h e e l 
 
 T h e   H L S   C o l o r   W h e e l   i s   a   m a p p i n g   o f   t h e   h u e   a n d   s a t u r a t i o n   c o m p o n e n t s   o f   a   c o l o r   f o r   a   g i v e n   l i g h t n e s s   v a l u e .   I t   i s   t h e   v i e w   l o o k i n g   d i r e c t l y   d o w n   a   c o n e   r e p r e s e n t i n g   t h e   H L S   c o l o r   m o d e l . 
 
 H u e   i s   m e a s u r e d   i n   i n c r e a s i n g   v a l u e s   a s   y o u   m o v e   c o u n t e r c l o c k w i s e   a r o u n d   t h e   C o l o r   W h e e l .   Z e r o ,   o r   r e d ,   i s   l o c a t e d   o n   t h e   r i g h t   s i d e   o f   t h e   C o l o r   W h e e l . 
 
 L i g h t n e s s   i s   s p e c i f i e d   w i t h   t h e   L i g h t n e s s   S l i d e r   B a r . 
 
 S a t u r a t i o n   i s   m e a s u r e d   f r o m   t h e   c e n t e r   o f   t h e   C o l o r   W h e e l   t o   t h e   p e r i m e t e r .   Z e r o   s a t u r a t i o n   i s   l o c a t e d   a t   t h e   c e n t e r . 
 
 
 T o   s p e c i f y   a   c o l o r   u s i n g   t h e   H L S   C o l o r   W h e e l : 
 
 1 .   S e l e c t   t h e   l i g h t n e s s   v a l u e   f o r   y o u r   c o l o r   b y   d r a g g i n g   t h e   i n d i c a t o r   o n   t h e   L i g h t   s l i d e r   b a r   o r   b y   t y p i n g   a   v a l u e   i n   t h e   p e r c e n t a g e   f i e l d . 
 
 A   l i g h t n e s s   v a l u e   o f   z e r o   r e p r e s e n t s   b l a c k ;   1 0 0   r e p r e s e n t s   w h i t e . 
 
 2 .   C l i c k   a n y w h e r e   i n   t h e   C o l o r   W h e e l   t o   c h o o s e   t h e   h u e   a n d   s a t u r a t i o n   m i x   o f   t h e   n e w   c o l o r . 
 
 T h e   c r o s s h a i r   t r a c k s   y o u r   s e l e c t i o n   i n   t h e   C o l o r   W h e e l .   T h e   i n d i c a t o r s   f o r   t h e   s l i d e r s   r e p r e s e n t i n g   t h e   h u e   a n d   s a t u r a t i o n   c o m p o n e n t s   m o v e   t o   r e f l e c t   y o u r   s e l e c t i o n . 
 
 T h e   C o l o r   B o x   a l s o   c h a n g e s   t o   r e f l e c t   y o u r   s e l e c t i o n .   
 
 
 
 N O T E S :   Y o u   c a n   a l s o   s p e c i f y   c o l o r s   d i r e c t l y   f r o m   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s . 
 
 Y o u   c a n   d e f i n e   d i t h e r i n g   f o r   a   c o l o r   b y   s e l e c t i n g   D e f a u l t   C o l o r   T o l e r a n c e s   f r o m   t h e   O p t i o n s   M e n u   o r   b y   s e l e c t i n g   t h e   C o l o r   T o l e r a n c e s   V i e w   f r o m   t h e   V i e w s   M e n u . 
 
 T o l e r a n c e s V i e w���� �L� O �  O p t i o n s M e n u
>�    �P  ����������  T o l e r a n c e s    
?#    \ O p t i o n s M e n u
?N   � V i e w s M e n u
?r 
  �  \\>>������"bu �X  `   C o l o r M o d e l s��
?�    �
N� " H� T h e   R G B / C M Y   C o l o r   P l a n e 
 
 T h e   C o l o r   P l a n e   i s   u s e d   t o   s e l e c t   a   c o l o r   u s i n g   t h e   R G B   o r   C M Y   c o l o r   m o d e l   a s   r e p r e s e n t e d   b y   a   c o l o r   c u b e . 
 
 T h e   C o l o r   P l a n e   i s   a   m a p p i n g   o f   t w o   p r i m a r y   c o l o r   c o m p o n e n t s   o f   a   c o l o r   f o r   a   g i v e n   v a l u e   o f   t h e   t h i r d   p r i m a r y   c o l o r   c o m p o n e n t .   I t   i s   a   v i e w   l o o k i n g   d i r e c t l y   d o w n   t h e   t o p   o f   t h e   c u b e   a t   a   p l a n e   d e t e r m i n e d   b y   t h e   v a l u e   o f   t h e   t h i r d   c o l o r   c o m p o n e n t . 
 
 T h e   c u b e   r e p r e s e n t s   e i t h e r   t h e   R G B   c o l o r   m o d e l   o r   t h e   C M Y   c o l o r   m o d e l . 
 
 I n   t h e   R G B   m o d e l ,   b y   d e f a u l t ,   t h e   g r e e n   a n d   b l u e   c o m p o n e n t s   a r e   m a p p e d   a g a i n s t   t h e   r e d   c o m p o n e n t .   I n   t h e   C M Y   m o d e l ,   t h e   m a g e n t a   a n d   y e l l o w   c o m p o n e n t s   a r e   m a p p e d   a g a i n s t   t h e   c y a n   c o m p o n e n t . 
 
 Y o u   c a n   c h a n g e   t h e   p l a n e   s e l e c t e d   f o r   v i e w i n g   t o   r e f l e c t   t h e   m a p p i n g   o f   a n y   t w o   p r i m a r y   c o l o r s   a g a i n s t   a   t h i r d   p r i m a r y   c o l o r .   U s e   t h e   c o l o r   p l a n e   o p t i o n s   i n   t h e   O p t i o n s   M e n u   t o   c h a n g e   t h e   d e f a u l t   m a p p i n g   o f   t h e   C o l o r   P l a n e . 
 
 T o   s p e c i f y   a   c o l o r   u s i n g   t h e   R G B   o r   C M Y   C o l o r   P l a n e : 
 
 1 .   C l i c k   a n y w h e r e   i n   t h e   C o l o r   P l a n e   t o   c h o o s e   a   v a l u e   f o r   t h e   t w o   c o l o r s   m a p p e d   i n   t h e   C o l o r   P l a n e . 
 
 T h e   c r o s s h a i r   t r a c k s   y o u r   s e l e c t i o n   a s   y o u   d r a g   t h e   p o i n t e r   i n   t h e   C o l o r   P l a n e .   T h e   i n d i c a t o r s   f o r   t h e   s l i d e r s   ( r e p r e s e n t i n g   t h e   t w o   m a p p e d   c o l o r s )   m o v e   t o   r e f l e c t   y o u r   s e l e c t i o n .   T h e   C o l o r   B o x   a l s o   c h a n g e s   t o   r e f l e c t   t h e   s e l e c t i o n . 
 
 2 .   M o v e   t h e   s l i d e r   f o r   t h e   t h i r d   c o m p o n e n t   t o   c h a n g e   i t s   v a l u e . 
 
 T h e   C o l o r   P l a n e   c h a n g e s   a s   y o u   m o v e   t h e   s l i d e r . 
 
 
 N O T E S :   Y o u   c a n   a l s o   s p e c i f y   c o l o r s   d i r e c t l y   f r o m   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s . 
 
 Y o u   c a n   d e f i n e   d i t h e r i n g   f o r   a   c o l o r   b y   s e l e c t i n g   D e f a u l t   C o l o r   T o l e r a n c e s   f r o m   t h e   O p t i o n s   M e n u   o r   b y   s e l e c t i n g   t h e   C o l o r   T o l e r a n c e s   V i e w   f r o m   t h e   V i e w s   M e n u . 
 
 
I N a m e d   C o l o r s 
 
 T h e   C o l o r   C h o o s e r   c o n t a i n s   a   s e t   o f   p r e d e f i n e d   c o l o r s   a v a i l a b l e   f o r   y o u r   u s e . 
 
 T h e s e   p r e d e f i n e d   c o l o r s   c a n   b e   s e l e c t e d   f r o m   t h e   c o l o r   l i s t   i n   t h e   N a m e d   C o l o r s   v i e w . 
 
 T h e   c o l o r s   i n   t h e   l i s t   c a n   b e   s o r t e d   b y   n a m e   o r   h u e   b y   s e l e c t i n g   t h e   a p p r o p r i a t e   o p t i o n   i n   t h e   O p t i o n s   M e n u . 
 
 
 R e f o r m S l i d e r s � C o n f i r m a t i o n   B u t t o n s 
 
 U s e   t h e   c o n f i r m a t i o n   b u t t o n s   t o   a p p l y   y o u r   s e l e c t i o n . 
 
��������� ����    C C c&a     �d  � C o l o r   T o l e r a n c e s   V i e w 
 
 U s e   t h e   C o l o r   T o l e r a n c e s   V i e w   t o   p r o v i d e   a d d e d   p r e c i s i o n   i n   d e f i n i n g   c o l o r   t o l e r a n c e s . 
 
 I n   t h e   C o l o r   T o l e r a n c e s   V i e w ,   u s e   t h e   D i t h e r   A r e a   o p t i o n   m e n u   t o   s e l e c t   a   d i t h e r i n g   m a t r i x .   U s e   t h e   D e l t a   V a l u e s   s l i d e r s   t o   s p e c i f y   a   d e l t a   v a l u e   f o r   e a c h   c o m p o n e n t   i n d i v i d u a l l y .   U s e   t h e   D i s t a n c e   s l i d e r   t o   s p e c i f y   a   d e l t a   v a l u e ,   o r   d i s t a n c e ,   t o   a p p l y   e q u a l l y   t o   a l l   c o m p o n e n t s . 
 
 F o r   m o s t   a p p l i c a t i o n s ,   t h e   c o l o r   t o l e r a n c e s   a v a i l a b l e   i n   t h e   D e f a u l t   C o l o r   T o l e r a n c e s   M e n u   ( i n   t h e   O p t i o n s   M e n u )   a r e   s u f f i c i e n t   t o   d e f i n e   y o u r   c o l o r s .   H o w e v e r ,   i f   y o u   r e q u i r e   m o r e   p r e c i s i o n   i n   d e f i n i n g   a   c o l o r ,   u s e   t h e   C o l o r   T o l e r a n c e s   V i e w   f r o m   t h e   V i e w s   M e n u .   
 
 C A U T I O N :   W h e n   s e l e c t i n g   a   d i t h e r i n g   m a t r i x ,   b e   c a r e f u l   a b o u t   s p e c i f y i n g   n o   d i t h e r i n g   f o r   a   c o l o r .   O n   m o s t   d i s p l a y s ,   s e l e c t i n g   t o o   m a n y   u n d i t h e r e d   c o l o r s   l i m i t s   t h e   n u m b e r   o f   c o l o r s   a v a i l a b l e   f o r   o t h e r   u s e s . 
 
 
8  H L S M o d e l��8�
V�    w"b� R G B M o d e l
V�   ; C M Y M o d e l
W   C G r a y s c a l e M o d e l
W4 	  :  ������	CC������	      �l  "?�� T o l e r a n c e s
W�   �	 ZZ__nn1e&���� �t  
]   
]$   <"?SE C o l o r   C o m p o n e n t   S l i d e r   B a r s 
 
 U s e   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s   t o   s p e c i f y   v a l u e s   f o r   i n d i v i d u a l   c o m p o n e n t s   o f   a   c o l o r .   
 
 T h e   c o l o r   c o m p o n e n t s   r e p r e s e n t e d   b y   t h e   s l i d e r   b a r s   v a r i e s   w i t h   e a c h   c o l o r   m o d e l .   E a c h   s l i d e r   b a r   h a s   a n   i n d i c a t o r   t h a t   d e f i n e s   t h e   v a l u e   o f   a   c o l o r   c o m p o n e n t . 
 
 T o   s p e c i f y   a   v a l u e   w i t h   a   s l i d e r   b a r ,   d o   o n e   o f   t h e   f o l l o w i n g : 
 
 * 	 D r a g   t h e   i n d i c a t o r   t o   t h e   d e s i r e d   l o c a t i o n   o n   t h e   s l i d e r 
 
 * 	 E n t e r   t h e   v a l u e   d i r e c t l y   i n t o   t h e   p e r c e n t a g e   f i e l d   f o r   t h e   s l i d e r 
 
 * 	 C l i c k   a n   a r e a   i n   t h e   s l i d e r   t o   s e l e c t   a   n e w   v a l u e 
 
 
 S e l e c t   R e f o r m   S l i d e r   I m a g e s   f r o m   t h e   O p t i o n s   M e n u   t o   d e f i n e   t h e   a p p e a r a n c e   a n d   b e h a v i o r   o f   t h e   s l i d e r   b a r s . 
 
 C o l o r W h e e l��8� C o l o r S l i d e r s	 kkpp{{1e�"Otg ���� �|  �� 1ef C o l o r P l a n e
]w   4 C o l o r S l i d e r s
]�   \	 nntt��
]�   <����   �  �       {{ C o l o r P l a n ed C o l o r S l i d e r s
^   d�����1������   �  �    !
^z   0���� O p t i o n s M e n u T o l e r a n c e s V i e w
^�   J V i e w s M e n u
^� 
  i" T o l e r a n c e s D e t a i l
^�   �
  �    "  FF`����BB  1eU%� i c �  �       �    ,  �    � �     b �   � � x     ;� �I �K{ �            W h e n   R e f o r m   S l i d e r   I m a g e s   i s   s e l e c t e d ,   t h e   s l i d e r   b a r s   d y n a m i c a l l y   r e f l e c t   t h e   a p p e a r a n c e   o f   t h e   c o l o r   b e i n g   s e l e c t e d .   A s   y o u   d r a g   t h e   i n d i c a t o r   t o   a   n e w   p o s i t i o n   o n   a n y   s l i d e r ,   t h e   a p p e a r a n c e   o f   t h e   o t h e r   s l i d e r s   c h a n g e s   t o   r e f l e c t   y o u r   s e l e c t i o n . 
 
 W h e n   R e f o r m   S l i d e r   I m a g e s   i s   n o t   s e l e c t e d ,   t h e   s l i d e r   b a r s   r e p r e s e n t   a n   u n c h a n g i n g   s c a l e   o f   v a l u e s   f o r   e a c h   c o m p o n e n t   o f   t h e   c o l o r . 
 
 � a-a!qaa
!aaaaqa	
!qqaaq!qaa!qa!aa !&!aaaa(!a,aaKqa9                                                         C o l o r   M o d e l s 
 
 F o u r   c o l o r   m o d e l s   a r e   a v a i l a b l e   f o r   c h o o s i n g   c o l o r s : 
 
 * 	 H L S 
 * 	 R G B 
 * 	 C M Y 
 * 	 G r a y s c a l e 
 
 H L S   C o l o r   M o d e l 
 T h e   H L S   c o l o r   m o d e l   s p e c i f i e s   a   c o l o r   u s i n g   a   c o m b i n a t i o n   o f   t h e   c o l o r ' s   h u e ,   l i g h t n e s s ,   a n d   s a t u r a t i o n   c o m p o n e n t s .   H L S   i s   t h e   d e f a u l t   c o l o r   m o d e l   f o r   t h e   C o l o r   C h o o s e r . 
 
 R G B   a n d   C M Y   C o l o r   M o d e l s 
 T h e   R G B   a n d   C M Y   c o l o r   m o d e l s   d e f i n e   c o l o r s   b y   s p e c i f y i n g   a   m i x t u r e   o f   p r i m a r y   c o l o r s . 
 
 T h e   R G B   m o d e l   m i x e s   t h e   a d d i t i v e   p r i m a r y   c o l o r s :   r e d ,   g r e e n ,   a n d   b l u e . 
 
 T h e   C M Y   m o d e l   m i x e s   t h e   s u b t r a c t i v e   p r i m a r y   c o l o r s :   c y a n ,   m a g e n t a ,   a n d   y e l l o w . 
 
 G r a y s c a l e   M o d e l 
 T h e   G r a y s c a l e   m o d e l   d e f i n e s   s h a d e s   o f   g r a y   f o r   b l a c k   a n d   w h i t e   o r   m o n o c h r o m e   m o n i t o r s . 
 
 � aaaq	AttributeContextaqBlock!untaQsExtraaKeywordBlockqLengthqasinkListqATypea	NodeBlockADataA	Texts!OffsetaasTag!extAAttributes	itleQsa
ypeVersionavhelpDocument�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                a G r a y s c a l e   C o l o r   M o d e l 
 
 T h e   G r a y s c a l e   m o d e l   d e f i n e s   s h a d e s   o f   g r a y   f o r   b l a c k   a n d   w h i t e   o r   m o n o c h r o m e   m o n i t o r s . 
 
 A   v a l u e   o f   1 0 0   i n   t h e   G r a y s c a l e   m o d e l   r e p r e s e n t s   w h i t e ;   z e r o   r e p r e s e n t s   b l a c k . 
 
 T h e   G r a y s c a l e   m o d e l   c a n   b e   r e p r e s e n t e d   a s   t h e   d i a g o n a l   l i n e   d r a w n   i n   t h e   R G B   c u b e   w h e n   t h e   v a l u e s   f o r   r e d ,   g r e e n ,   a n d   b l u e   a r e   e q u a l . 
 
 T h e   G r a y s c a l e   s l i d e r   b a r   c o r r e s p o n d s   t o   t h i s   d i a g o n a l   l i n e . 
 
 T o   s p e c i f y   a   c o l o r   i n   t h e   G r a y s c a l e   M o d e l ,   d o   a n y   o f   t h e   f o l l o w i n g : 
 
 * 	 D r a g   t h e   i n d i c a t o r   t o   t h e   d e s i r e d   v a l u e   o f   t h e   G r a y s c a l e   s l i d e r . 
 
 * 	 C l i c k   o n   t h e   d e s i r e d   v a l u e   i n   t h e   G r a y s c a l e   s l i d e r . 
 
 * 	 S p e c i f y   a   v a l u e   i n   t h e   p e r c e n t a g e   f i e l d   o f   t h e   G r a y s c a l e   s l i d e r . 
 
 
 I n   a l l   i n s t a n c e s ,   t h e   C o l o r   B o x   c h a n g e s   t o   r e f l e c t   y o u r   s e l e c t i o n . 
 
 N O T E S :   T h e   C o l o r   V i e w   a r e a   i s   i n a c t i v e   w h e n   s p e c i f y i n g   c o l o r s   w i t h   t h e   G r a y s c a l e   M o d e l . 
 
 I f   t h e   C o l o r   B o x   d i s p l a y s   y o u r   s e l e c t i o n s   o n l y   a s   s o l i d   b l a c k   o r   s o l i d   w h i t e ,   y o u   m a y   h a v e   t o   s p e c i f y   c o l o r   t o l e r a n c e s   f o r   d i t h e r i n g . 
 
 
 
 
 �                                                                                                                                                           � H L S   C o l o r   M o d e l 
 
 T h e   H L S   c o l o r   m o d e l   d e f i n e s   a   c o l o r   b y   s p e c i f y i n g   v a l u e s   f o r   t h e   c o l o r ' s   h u e ,   l i g h t n e s s ,   a n d   s a t u r a t i o n   c o m p o n e n t s .   T h e s e   c o m p o n e n t s   c a n   b e   r e p r e s e n t e d   a s   a   " c o l o r   c o n e . " 
 
 T h e   h u e   c o m p o n e n t   d e f i n e s   a   c o l o r ' s   p o s i t i o n   i n   a   c o n t i n u o u s   c o l o r   s p e c t r u m ,   a n d   i s   r e p r e s e n t e d   a s   t h e   a n g l e   a r o u n d   t h e   c i r c u m f e r e n c e   o f   t h e   c o n e .   H u e   i s   m e a s u r e d   i n   d e g r e e s   a n d   r a n g e s   f r o m   z e r o   t o   3 6 0 .   Z e r o   r e p r e s e n t s   r e d . 
 
 T h e   l i g h t n e s s   c o m p o n e n t   d e f i n e s   t h e   d e n s i t y   o f   a   c o l o r   a n d   i s   r e p r e s e n t e d   b y   t h e   v e r t i c a l   a x i s   o f   t h e   c o n e .   L i g h t n e s s   r a n g e s   f r o m   z e r o   f o r   b l a c k ,   t o   1 0 0   f o r   w h i t e . 
 
 S a t u r a t i o n   d e f i n e s   t h e   i n t e n s i t y   o f   a   c o l o r   a n d   i s   r e p r e s e n t e d   b y   t h e   d i s t a n c e   f r o m   t h e   v e r t i c a l   a x i s   t o   t h e   p e r i m e t e r   o f   t h e   c o n e .   S a t u r a t i o n   r a n g e s   f r o m   z e r o   t o   1 0 0 . 
 
 T o   s p e c i f y   a   c o l o r   i n   t h e   H L S   M o d e l   u s e   t h e   C o l o r   W h e e l   i n   c o m b i n a t i o n   w i t h   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s . 
 
G                                                                                                                                                                                                                                                                                                                                     � R G B   C o l o r   M o d e l 
 
 T h e   R G B   c o l o r   m o d e l   d e f i n e s   c o l o r s   b y   s p e c i f y i n g   a   m i x t u r e   o f   t h e   a d d i t i v e   p r i m a r y   c o l o r s   r e d ,   g r e e n ,   a n d   b l u e . 
 
 T h e   R G B   c o l o r   m o d e l   c a n   b e   r e p r e s e n t e d   a s   a   " c o l o r   c u b e . "   T h e   h e i g h t ,   w i d t h ,   a n d   l e n g t h   o f   t h e   c u b e   e a c h   r e p r e s e n t   a   p r i m a r y   c o l o r . 
 
 T o   s p e c i f y   a   c o l o r   i n   t h e   R G B   M o d e l ,   u s e   t h e   R G B   C o l o r   P l a n e   i n   c o m b i n a t i o n   w i t h   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s . 
 
 
 
 
                                                                                                                                                                                                                                                                C M Y   C o l o r   M o d e l 
 
 T h e   C M Y   c o l o r   m o d e l   d e f i n e s   c o l o r s   b y   s p e c i f y i n g   a   m i x t u r e   o f   t h e   s u b t r a c t i v e   p r i m a r y   c o l o r s   c y a n ,   m a g e n t a ,   a n d   y e l l o w . 
 
 T h e   C M Y   c o l o r   m o d e l   c a n   b e   r e p r e s e n t e d   a s   a   " c o l o r   c u b e . "   T h e   h e i g h t ,   w i d t h ,   a n d   l e n g t h   o f   t h e   c u b e   e a c h   r e p r e s e n t   a   p r i m a r y   c o l o r . 
 
 T o   s p e c i f y   a   c o l o r   i n   t h e   C M Y   M o d e l ,   u s e   t h e   C M Y   C o l o r   P l a n e   i n   c o m b i n a t i o n   w i t h   t h e   C o l o r   C o m p o n e n t   S l i d e r   B a r s . 
 
 
 
 
 �                                                                                                                                                                                                                                               � C o l o r   T o l e r a n c e s 
 
 S i n c e   m a n y   d i s p l a y s   c a n n o t   a c c u r a t e l y   r e p r e s e n t   a l l   c o l o r s ,   d i t h e r i n g   i s   u s e d   t o   a p p r o x i m a t e   c o l o r s   o n   a   d i s p l a y .   D i t h e r i n g   t a k e s   p l a c e   w i t h i n   c e r t a i n   t o l e r a n c e s   y o u   d e f i n e   i n   t h e   C o l o r   C h o o s e r . 
 
 S p e c i f y   t h e   t o l e r a n c e s   f o r   d i t h e r i n g   c o l o r s   f r o m   t h e   D e f a u l t   C o l o r   T o l e r a n c e s   M e n u   i n   t h e   O p t i o n s   M e n u ,   o r   f r o m   t h e   C o l o r   T o l e r a n c e s   V i e w   f r o m   t h e   V i e w s   M e n u . 
 
 F o r   m o s t   a p p l i c a t i o n s ,   t h e   d e f a u l t   v a l u e s   f o r   c o l o r   t o l e r a n c e s   a v a i l a b l e   i n   t h e   D e f a u l t   C o l o r   T o l e r a n c e s   M e n u   a r e   s u f f i c i e n t   t o   d e f i n e   y o u r   c o l o r s .   H o w e v e r ,   i f   y o u   r e q u i r e   m o r e   p r e c i s i o n   i n   d e f i n i n g   a   c o l o r ,   u s e   t h e   C o l o r   T o l e r a n c e s   V i e w   f r o m   t h e   V i e w s   M e n u .   
 
 C A U T I O N :   W h e n   s e l e c t i n g   a   d i t h e r i n g   m a t r i x ,   b e   c a r e f u l   a b o u t   s p e c i f y i n g   n o   d i t h e r i n g   f o r   a   c o l o r .   O n   m o s t   d i s p l a y s ,   s e l e c t i n g   t o o   m a n y   c o l o r s   t h a t   a r e   n o t   d i t h e r e d   l i m i t s   t h e   n u m b e r   o f   c o l o r s   a v a i l a b l e   f o r   o t h e r   u s e s . 
 
 
 
 
I                                                                                                                                                                                                                                                                                                                                       � D e f a u l t   C o l o r   T o l e r a n c e s   D e t a i l s 
 
 T h e   s e l e c t i o n s   a v a i l a b l e   f r o m   t h e   D e f a u l t   C o l o r   T o l e r a n c e s   m e n u   p r o v i d e   t h e   p r e c i s i o n   n e e d e d   i n   m o s t   a p p l i c a t i o n s .   T h e   c o l o r   t o l e r a n c e   v a l u e s   c o r r e s p o n d i n g   t o   t h e s e   m e n u   s e l e c t i o n s   a r e   l i s t e d   b e l o w .   T h e   s i z e   o f   t h e   d i t h e r   a r e a   a n d   d i t h e r i n g   p e r c e n t a g e   i s   l i s t e d   b e n e a t h   e a c h   s p e c i f i c a t i o n .   
 
 D e f a u l t   C o l o r   T o l e r a n c e s 
 
 L a r g e   D i t h e r 
 8   x   8   
 . 3 9   p e r c e n t 
 
 S m a l l   D i t h e r 
 2   x   2 
 6 . 2 5   p e r c e n t 
 
 S o l i d 
 N o   D i t h e r i n g 
 2 5 . 0 0   p e r c e n t 
 
 P r e c i s e   L a r g e   D i t h e r 
 1 6   x   1 6 
 0 . 1 9   p e r c e n t 
 
 P r e c i s e   S m a l l   D i t h e r 
 4   x   4 
 1 . 5 6   p e r c e n t 
 
 P r e c i s e   S o l i d 
 N o   D i t h e r i n g 
 6 . 2 5   p e r c e n t 
 
 
 C A U T I O N :   B e   c a r e f u l   w h e n   s e l e c t i n g   S o l i d   o r   P r e c i s e   S o l i d   f r o m   t h e   C o l o r   T o l e r a n c e s   m e n u .   T h e s e   s e l e c t i o n s   s p e c i f y   t h a t   n o   d i t h e r i n g   t a k e   p l a c e .   O n   m o s t   d i s p l a y s ,   s e l e c t i n g   t o o   m a n y   u n d i t h e r e d   c o l o r s   l i m i t s   t h e   n u m b e r   o f   c o l o r s   a v a i l a b l e   f o r   o t h e r   u s e s . 
 
y                                                                                                                                                                                                                                                                                                                                                                                       w�� �ab b�AabNR �r
�b�bZbPaa"KaqGbx"(jb&3�b&?7r&I�r&VMB&\jr&h�B&q"�r&{#b& �b#�&b �>�b& �r?&r �?�b>�r&O�r& �bO�&b �Wy"& �bW�&b �]Vb& �b]�&" �^Nr& �b^p&ab�!#!!R#Ua#a%b#�b�b,(�",(
�r,(	b,(-b,(Mb,(ub,(�",(�r,(�b,(�r(�b,(�b�r�bsb�b3�",9	",9Mb,9s",9�",9�b(?b,9+"�" b�b�b?0b,Enb,E�",E�r(eb,E�b�b"8bBbISb,Oz,O�b,O�r,O�b,OR,OBr�b,O�Bb�rH�"(r"UrbbfYb\{b,a�r,a�r,a2,a+",aSb,ay(�b,a�B�b�r��2h�b,n�b,n"�R("�b,n"�B]b"�r"��rq"�,w#2,w#[r,w#�r(#�r,w#7r#�b#�"#�b#�2{#�2, �"#�," �&�r, �b&�, �&�b('b, �b&}a&�!B#�ab'ab'" �'", �r':,b �'|, �B'�,B �'�2, �b'�,b �'�b(>�r, �b'Xab�qb'�!R'�ab'r ��r, �b>�(!R?ab�qb>�qb'"Ab>�r �?b, �r?C,b �?�"(?�r, �R?gqb?�ab?�qb?�q"?:b �?b, �r?�q"?�," �?�r?b?�rO�"?�b(O�BO�bO�bO�bO�" �bO�,b �V�b, �rW)," �WSb(W�b, �rWqbW^abWoqrV�abW�r �O�b, �bW�(abW�abW�abW�q"W�abV�b �V�", �rW�(qb]^," �W�b]?qW�]IV� �], �]�(]�, �]� ]� ]N ]r ]  �]g, �]�(^V, �^1!]�!^!^G!]l �^<, �^e, �^�, �_ _, �^�"_"_/"_B"_= �