��     4  {�d  �sw    I m a g e   E d i t o r F i l e   M e n u"� I m a g e   E d i t o r& I m a g e   E d i t i n g   A r e a  ��� ��  ��   ��   ��   ��   ��   ��     	 ����  �� 
  ��      ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ����     ����  ��    �� ��   �� ! �� " �� # �� $ ���� I m a g e   F o r m a t sL ^� y�"a E����'H]x���� $9Tq���,K~���,4 T r a n s p a r e n c y   E d i t i n g   A r e a> I m p o r t i n g   a n d   E x p o r t i n g   I m a g e s, S e t   I m a g e   S i z e   W i n d o w E d i t   M e n u8 S e l e c t i n g   A r e a s   f o r   E d i t i n g V i e w   M e n u O p t i o n s   M e n u T o o l   P a l e t t e  K e y b o a r d   M a c r o s H a n d   T o o l D r o p p e r   T o o l S e l e c t i o n   T o o l L a s s o   T o o l F i l l   T o o l S p r a y   C a n   T o o l E r a s e r   T o o l4  T e x t   T o o l P e n c i l L i n e   T o o l E l l i p s e   T o o l S o l i d   E l l i p s e R e c t a n g l e   T o o l  S o l i d   R e c t a n g l e C o l o r   P a l e t t e6 S e t t i n g   C o l o r s   f o r   D r a w i n g& L i n e   W i d t h   P a l e t t e P a l e t t e   E d i t o r2 P a l e t t e   E d i t o r   F i l e   M e n u2 P a l e t t e   E d i t o r   E d i t   M e n u P a l e t t e s   M e n u, C o l o r   P a l e t t e   B u t t o n s0 E d i t i n g   a   C o l o r   P a l e t t e6 I n s t a l l i n g   a   C o l o r   P a l e t t e��
�
�  P e n c i l ' E d i t M e n uP�_x��p���� !6Wf�������		-	L	a	|	�	�	�	�


C
^
q
� O v e r v i e w  I m a g e E d i t o r L i n e W i d t h P a l)  "!
$#	  T o o l P a l e t t e S e t t i n g C o l o r s C o l o r P a l e t t e H a n d T o o l R e c t T o o l L i n e T o o l E r a s e r%   C o l o r P a l B u t t o n s S p r a y T o o l  C o l o r P a l P a l M e n u P a l e E d" I m p o r t E x p o r t P r o c S o l R e c t S i z e W i n d o w S o l E l l i p s e T e x t T o o l F i l e M e n u M a c r o s O p t i o n s M e n u S e l e c t A r e a T r a n s p E d i t A r e a L a s s o T o o l I m a g e F o r m a t s I m a g e E d i t A r e a D r o p T o o l" C o l o r P a l F i l e M e n u F i l l T o o l  I n s t a l l C o l o r P a l S e l T o o l. I m a g e E d i t o r P a l e d D i a l o g E d i t C o l o r P a l V i e w M e n u E l l i p s e" C o l o r P a l E d i t M e n u    *   p a l e t t e   e d i t o r i m a g e   e d i t o r
G   5643
k 	   �   7  28G9:;<=>?@ABCDE�  I m a g e F o r m a t s
M   H" I m p o r t E x p o r t P r o c
s    e F i l e M e n u
� 	   � E d i t M e n u
� 	   � V i e w M e n u
� 	   �I = I m a g e   E d i t o r 
 
 U s e   t h e   I m a g e   E d i t o r   t o   c r e a t e   a n d   e d i t   i m a g e s   i n   v a r i o u s   i m a g e   f o r m a t s . 
 
 Y o u   c a n   a l s o   i m p o r t   a n d   e x p o r t   i m a g e s   t o   a n d   f r o m   t h e   I m a g e   E d i t o r . 
 
 T h e   f o l l o w i n g   c o m p o n e n t s   a r e   v i s i b l e   w h e n   t h e   I m a g e   E d i t o r   f i r s t   o p e n s : 
 
 F i l e   M e n u 
 E d i t   M e n u 
 V i e w   M e n u 
 O p t i o n s   M e n u 
 T o o l   P a l e t t e 
 C o l o r   P a l e t t e 
 I m a g e   E d i t i n g   A r e a 
 L i n e   W i d t h   P a l e t t e 
 F o r e g r o u n d   C o l o r   S e l e c t i o n   B o x 
 B a c k g r o u n d   C o l o r   S e l e c t i o n   B o x 
 
 T h e   f o l l o w i n g   c o m p o n e n t s   a r e   a v a i l a b l e   w h i l e   u s i n g   t h e   I m a g e   E d i t o r : 
 
 S e t   I m a g e   S i z e   W i n d o w 
 C o l o r   P a l e t t e   E d i t o r 
 T r a n s p a r e n c y   E d i t i n g   A r e a 
 
8MO O p t i o n s M e n uH  T o o l P a l e t t e
i    C o l o r P a l e t t e
�    I m a g e E d i t A r e a
�   , L i n e W i d t h P a l
�   ? C o l o r P a l e t t e
   R C o l o r P a l e t t e
'   q S i z e W i n d o w
M   � P a l e E d
o   � T r a n s p E d i t A r e a
�   % T h e   I m a g e   E d i t o r   s u p p o r t s   t h e   f o l l o w i n g   i m a g e   f o r m a t s : 
 
 
 B M P 	 P B M 
 
 D I B 	 P G M 
 
 G I F 	 P P M 
 
 I C O 	 X B M 
 
 
 R u n - l e n g t h   e n c o d e d   D I B   f o r m a t s   a r e   n o t   s u p p o r t e d .   
 L  8 JKIH
� 	   � T o o l P a l e t t e
' 	  01e&U  V i e w M e n u(     1 1;;	&&RSQP T  \^eX T o o l P a l e t t e
}   �      ��YZXW [$  
�   � I m a g e F o r m a t s
�  X ^^{ I m a g e   E d i t i n g   A r e a 
 
 T h e   I m a g e   E d i t i n g   A r e a   d i s p l a y s   t h e   i m a g e   c u r r e n t l y   b e i n g   e d i t e d .   I f   t h e   i m a g e   i s   t o o   l a r g e   t o   d i s p l a y   c o m p l e t e l y ,   y o u   c a n   u s e   t h e   s c r o l l   b a r s   o r   t h e   H a n d   T o o l   t o   s c r o l l   t h e   i m a g e . 
 
 V a r i o u s   o p t i o n s   d e f i n i n g   t h e   b e h a v i o r   a n d   a p p e a r a n c e   o f   t h e   I m a g e   E d i t i n g   A r e a   a r e   a v a i l a b l e   f r o m   t h e   V i e w   M e n u . 
 
,   I m a g e F o r m a t s1e   8  �o(ab`_ h0      : ���]"Yd�fgedilj I m a g e F o r m a t s
�  � I m a g e F o r m a t s
   S i z e W i n d o w
<   z   opnm��   : ? � � � � �*c�		 q<  	rystuvw S e l e c t A r e a *�
�   �(�� 
#�  
#�  F� T r a n s p a r e n c y   E d i t i n g   A r e a 
 
 S o m e   a p p l i c a t i o n s   u s e   t r a n s p a r e n c i e s   o f   i m a g e s   s o   t h a t   i m a g e s   a r e   d r a w n   p r o p e r l y   a g a i n s t   d i f f e r e n t   b a c k g r o u n d s .   T r a n s p a r e n c i e s   a r e   c r e a t e d   a n d   e d i t e d   i n   t h e   T r a n s p a r e n c y   E d i t i n g   A r e a . 
 
 W h e n   y o u   c r e a t e   a   t r a n s p a r e n c y   f o r   a n   i m a g e ,   y o u   c r e a t e   a   b l a c k   a n d   w h i t e   m a s k   f o r   t h e   i m a g e .   A r e a s   i n   t h e   o r i g i n a l   i m a g e   t h a t   a r e   n o t   b l a c k   a r e   m a s k e d   o u t   b y   t h e   b l a c k   a r e a   o f   t h e   t r a n s p a r e n c y .   T h i s   p r e v e n t s   b a c k g r o u n d   c o l o r s   f r o m   i n t e r f e r i n g   w i t h   y o u r   i m a g e .   T h e   w h i t e   a r e a s   o f   t h e   t r a n s p a r e n c y   a r e   c l e a r ,   a n d   d e f i n e   t h e   b l a c k   a r e a s   o f   t h e   o r i g i n a l   i m a g e . 
 
 T o   c r e a t e   a   t r a n s p a r e n c y   f o r   a n   i m a g e : 
 
 1 .   S e l e c t   C r e a t e   T r a n s p a r e n c y   f r o m   t h e   O p t i o n s   M e n u . 
 
 A   T r a n s p a r e n c y   E d i t i n g   A r e a   a p p e a r s . 
 
 2 .   U s i n g   t h e   S e l e c t i o n   T o o l s ,   s e l e c t   t h e   a r e a   o f   t h e   o r i g i n a l   i m a g e   y o u   w a n t   t o   m a s k . 
 
 D o u b l e - c l i c k   t h e   S e l e c t i o n   T o o l   t o   s e l e c t   t h e   e n t i r e   i m a g e . 
 
 3 .   S e l e c t   M a s k   S e l e c t i o n   f r o m   t h e   E d i t   M e n u . 
 
 A   m a s k   i s   c r e a t e d   f o r   t h e   s e l e c t e d   a r e a ,   a n d   d i s p l a y e d   i n   t h e   T r a n s p a r e n c y   E d i t i n g   A r e a .   T h i s   m a s k   i s   a   s t a r t i n g   p o i n t   f o r   c r e a t i n g   a   f i n a l   m a s k .   A n y   a r e a   o f   y o u r   i m a g e   c o n t a i n i n g   t h e   b a c k g r o u n d   c o l o r   i s   m a s k e d   o u t . 
 
 4 .   U s e   a n y   o f   t h e   t o o l s   f r o m   t h e   T o o l   P a l e t t e   t o   e d i t   t h e   t r a n s p a r e n c y ,   i f   n e c e s s a r y . 
 
 W h e n   e d i t i n g   a   t r a n s p a r e n c y ,   t h e   f o r e g r o u n d   c o l o r   i s   a l w a y s   s e t   t o   b l a c k   a n d   t h e   b a c k g r o u n d   c o l o r   t o   w h i t e . 
 
 
 T o   r e m o v e   a   t r a n s p a r e n c y : 
 
 1 .   S e l e c t   D e l e t e   T r a n s p a r e n c y   f r o m   t h e   O p t i o n s   M e n u . 
 
 T h e   T r a n s p a r e n c y   E d i t i n g   A r e a   i s   r e m o v e d   f r o m   t h e   I m a g e   E d i t o r   a n d   t h e   t r a n s p a r e n c y   i s   d e l e t e d . 
 
 S e l e c t A r e a S e l e c t A r e a S e l e c t A r e a
#�  } �D   5 I m p o r t i n g   a n d   E x p o r t i n g   I m a g e s 
 
 T o   i m p o r t   a n   i m a g e : 
 
 1 .   F r o m   t h e   F i l e   M e n u ,   s e l e c t   I m p o r t . . . 
 
 A   f i l e   c h o o s e r   a p p e a r s . 
 
 2 .   U s e   t h e   F i l t e r s   o p t i o n   i n   t h e   f i l e   c h o o s e r   t o   s p e c i f y   a n   i m a g e   f o r m a t . 
 
 T h e   f i l e   c h o o s e r   f i l t e r s   f i l e s   a c c o r d i n g   t o   y o u r   s p e c i f i c a t i o n . 
 
 3 .   S e l e c t   t h e   f i l e   y o u   w a n t   t o   i m p o r t ,   a n d   a p p l y   y o u r   s e l e c t i o n   i n   t h e   f i l e   c h o o s e r . 
 
 T h e   i m a g e   f r o m   t h e   t h e   f i l e   a p p e a r s   i n   t h e   I m a g e   E d i t o r . 
 
 
 T o   e x p o r t   a n   i m a g e : 
 
 1 .   F r o m   t h e   F i l e   M e n u ,   s e l e c t   E x p o r t . . . 
 
 A   f i l e   c h o o s e r   a p p e a r s . 
 
 2 .   I m a g e s   c a n   b e   e x p o r t e d   i n   v a r i o u s   i m a g e   f o r m a t s .   U s e   t h e   F i l t e r s   o p t i o n   i n   t h e   f i l e   c h o o s e r   t o   s p e c i f y   a n   i m a g e   f o r m a t   f o r   t h e   e x p o r t e d   f i l e . 
 
 3 .   S p e c i f y   t h e   p a t h   a n d   f i l e   n a m e   f o r   y o u r   e x p o r t e d   f i l e   i n   t h e   f i l e   c h o o s e r   a n d   a p p l y   y o u r   s e l e c t i o n . 
 
 T h e   i m a g e   i s   e x p o r t e d   t o   t h e   s e l e c t e d   d e s t i n a t i o n . 
 
 S e l e c t A r e a
*6  � T r a n s p E d i t A r e a
*X   � S e l e c t A r e a
*�  2 � U s e   t h e   S e l e c t i o n   T o o l   o r   L a s s o   T o o l   f r o m   t h e   T o o l   P a l e t t e   t o   s e l e c t   a r e a s   f o r   e d i t i n g .   
 T o o l P a l e t t e
+Z    .���~}|$$ &   :nnR�../Z���?���aa & 	   / / 	 ii         ���� S e t   I m a g e   S i z e   W i n d o w 
 
 T h e   S e t   I m a g e   S i z e   W i n d o w   s p e c i f i e s   t h e   s i z e   o f   a n   i m a g e   ( i n   p i x e l s ) . 
 
 T o   s p e c i f y   t h e   s i z e   o f   a n   i m a g e : 
 
 1 .   S e l e c t   S e t   S i z e   f r o m   t h e   F i l e   M e n u . 
 
 T h e   S e t   I m a g e   S i z e   W i n d o w   o p e n s . 
 
 2 .   S p e c i f y   t h e   w i d t h   a n d   h e i g h t   o f   t h e   i m a g e   i n   p i x e l s ,   a n d   s e l e c t   O K . 
 
 T h e   s i z e   o f   t h e   i m a g e   i n   t h e   I m a g e   E d i t o r   c h a n g e s   t o   r e f l e c t   y o u r   s e l e c t i o n ,   a n d   t h e   S e t   I m a g e   S i z e   W i n d o w   c l o s e s . 
               T o o l P a l e t t e
/#   ` T o o l P a l e t t e
/G 	  �   @ �<P �T   T o o l P a l e t t e 
/� 	   � P a l e E d
/�    �  oo T r a n s p E d i t A r e a
/�    � F i l e   M e n u 
 
 T h e   F i l e   M e n u   c o n t a i n s   t h e   f o l l o w i n g   o p t i o n s : 
 
 C l o s e 
 C l o s e s   t h e   I m a g e   E d i t o r .   T h e   i m a g e   c u r r e n t l y   b e i n g   e d i t e d   i s   a p p l i e d   i n   t h e   a p p l i c a t i o n . 
 
 S a v e 
 T h e   i m a g e   c u r r e n t l y   b e i n g   e d i t e d   i s   a p p l i e d   i n   t h e   a p p l i c a t i o n ,   b u t   t h e   I m a g e   E d i t o r   d o e s   n o t   c l o s e . 
 
 I m p o r t 
 I m p o r t s   a n   i m a g e .   W h e n   t h i s   o p t i o n   i s   s e l e c t e d   a   f i l e   c h o o s e r   o p e n s .   U s e   t h e   f i l e   c h o o s e r   t o   s e l e c t   a n   i m a g e   t o   i m p o r t .   
 
 T h e   F i l t e r s   o p t i o n   i n   t h e   f i l e   c h o o s e r   a l l o w s   y o u   t o   s e l e c t   a n   i m a g e   f o r m a t   t o   d i s p l a y   i n   t h e   f i l e   c h o o s e r . 
 
 E x p o r t 
 W r i t e s   t h e   c u r r e n t   i m a g e   t o   a   f i l e .   W h e n   t h i s   o p t i o n   i s   s e l e c t e d   a   f i l e   c h o o s e r   o p e n s .   U s e   t h e   f i l e   c h o o s e r   t o   s e l e c t   a   l o c a t i o n   a n d   i m a g e   f o r m a t   f o r   t h e   e x p o r t e d   f i l e . 
 
 S e t   S i z e . . . 
 U s e   t h i s   o p t i o n   t o   s p e c i f y   a   s i z e   f o r   a n   i m a g e . 
 
 W h e n   t h i s   o p t i o n   i s   s e l e c t e d ,   t h e   S e t   I m a g e   S i z e   W i n d o w   o p e n s .   S p e c i f y   a   s i z e   f o r   y o u r   i m a g e   i n   t h e   S e t   I m a g e   S i z e   W i n d o w . 
 
 R e v e r t 
 R e s t o r e s   t h e   I m a g e   E d i t o r   t o   t h e   l a s t   s a v e d   v e r s i o n .   A l l   c h a n g e s   m a d e   t o   t h e   e d i t o r   s i n c e   t h e   l a s t   s a v e d   v e r s i o n   a r e   l o s t . 
 
 N o t e   t h a t   t h e   c o n t e n t s   o f   t h e   I m a g e   E d i t o r   a r e   a l s o   c o n s i d e r e d   " s a v e d "   a f t e r   t h e   C l o s e   c o m m a n d   ( f r o m   t h e   F i l e   M e n u )   i s   i s s u e d . 
 
 
1% �\  �������������������� M a c r o sd  
8�    u H a n d T o o l
9   � D r o p T o o l
9/   � S e l T o o l
9M 	  � L a s s o T o o l
9i   � F i l l T o o l
9�   � S p r a y T o o l
9�   � E r a s e r
9�   � T e x t T o o l
9�   P e n c i l
9�   L i n e T o o l
:   E l l i p s e
:7    S o l E l l i p s e
:S  - R e c t T o o l
:u 	 E S o l R e c t
:�  S M a c r o s
:�   R  ��( e������ @� "	 � �����"���� �Y>  C o l o r P a l e t t ea 
;6    �� "B* ����B�  "
����� Q� � "	 �  ����i> "����� l   � " � p  !� E d i t   M e n u 
 
 T h e   E d i t   M e n u   c o n t a i n s   t h e   f o l l o w i n g   o p t i o n s : 
 
 U n d o 
 R e d o 
 U s e   t h e s e   o p t i o n s   t o   u n d o   o r   r e d o   e d i t i n g   a c t i o n s   i n   t h e   I m a g e   E d i t o r . 
 
 C u t 
 C o p y 
 P a s t e 
 C l e a r 
 U s e   t h e s e   o p t i o n s   t o   p e r f o r m   e d i t i n g   a c t i o n s   o n   s e l e c t e d   a r e a s   i n   t h e   I m a g e   E d i t i n g   A r e a . 
 
 R o t a t e 
 R o t a t e s   t h e   s e l e c t e d   a r e a   9 0   d e g r e e s . 
 
 F l i p   H o r i z o n t a l 
 M i r r o r s   t h e   s e l e c t e d   a r e a   h o r i z o n t a l l y . 
 
 F l i p   V e r t i c a l 
 M i r r o r s   t h e   s e l e c t e d   a r e a   v e r t i c a l l y . 
 
 M a s k   S e l e c t i o n 
 C r e a t e s   a   m a s k   o f   t h e   s e l e c t e d   a r e a . 
 T h i s   o p t i o n   i s   o n l y   a v a i l a b l e   w h e n   c r e a t i n g   a   t r a n s p a r e n c y . 
 
 C r o p   t o   S e l e c t i o n 
 C r o p s   t h e   i m a g e   t o   t h e   s e l e c t e d   a r e a . 
 
� H a n d   T o o l 
 
 U s e   t h e   H a n d   T o o l   t o   r e p o s i t i o n   t h e   v i s i b l e   p a r t   o f   t h e   i m a g e   w h e n   a n   o v e r s i z e   i m a g e   i s   i n   t h e   I m a g e   E d i t i n g   A r e a . 
 
 S e l e c t   a n d   d r a g   t h e   o v e r s i z e   i m a g e   w i t h   t h e   H a n d   T o o l   t o   r e p o s i t i o n   t h e   i m a g e .   
M L a s s o   T o o l 
 
 U s e   t h e   L a s s o   T o o l   t o   s e l e c t   a n y   i r r e g u l a r   a r e a   o f   a n   i m a g e   f o r   e d i t i n g . 
 
 D r a g   t h e   p o i n t e r   w i t h   t h e   L a s s o   T o o l   t o   s u r r o u n d   t h e   a r e a   y o u   w a n t   t o   s e l e c t .   
����� "	 �  ����t  ""&����� q� #� "	 �  ����x  $"����� � V i e w   M e n u 
 
 T h e   V i e w   M e n u   c o n t a i n s   t h e   f o l l o w i n g   o p t i o n s : 
 
 F a t   B i t s 
 M a g n i f i e s   t h e   i m a g e   i n   t h e   I m a g e   E d i t i n g   A r e a   s o   e a c h   p i x e l   c a n   b e   v i e w e d . 
 
 T h e   d e f a u l t   m a g n i f i c a t i o n   w h e n   F a t   B i t s   i s   e n a b l e d   i s   5 x .   W h e n   F a t   B i t s   i s   d i s a b l e d ,   t h e   i m a g e   r e t u r n s   t o   i t s   a c t u a l   s i z e . 
 
 D r a w   F r o m   C e n t e r 
 D e f i n e s   t h e   s t a r t i n g   p o i n t   f o r   t h e   f o l l o w i n g   d r a w i n g   t o o l s   f r o m   t h e   T o o l   P a l e t t e : 
 
 * 	 L i n e   T o o l 
 * 	 E l l i p s e   T o o l s 
 * 	 R e c t a n g l e   T o o l s 
 
 N o r m a l l y   t h e s e   t o o l s   b e g i n   d r a w i n g   a n   i t e m   f r o m   t h e   e n d   ( o r   p e r i m e t e r )   o f   t h e   i t e m .   S e l e c t i n g   t h e   D r a w   F r o m   C e n t e r   o p t i o n   s p e c i f i e s   t h a t   d r a w i n g   b e g i n s   a t   t h e   c e n t e r   o f   t h e   i t e m . 
 
 S h o w   G r i d 
 D i s p l a y   t h e   i m a g e   i n   a   g r i d .   I n d i v i d u a l   p i x e l s   a r e   o u t l i n e d   w i t h   t h e   g r i d   p a t t e r n .   W h e n   t h e   b i t   s i z e   i s   s m a l l e r   t h a n   t h r e e   p i x e l s ,   t h e   g r i d   i s   n o t   s h o w n . 
 
 S h o w   P o s i t i o n 
 D i s p l a y s   t h e   c o o r d i n a t e s   o f   a n   i m a g e   a b o v e   t h e   I m a g e   E d i t i n g   A r e a . 
 
 T h e   c o o r d i n a t e s   p r o v i d e   i n f o r m a t i o n   o n   t h e   p o s i t i o n ,   d i r e c t i o n ,   a n d   s i z e   o f   e d i t i n g   o p e r a t i o n s .   T h e   o r i g i n   o f   t h e   i m a g e   i s   t h e   l o w e r   l e f t   c o r n e r   o f   t h e   i m a g e . 
 
 T h e   f o l l o w i n g   i n f o r m a t i o n   i s   d i s p l a y e d   b y   t h e   S h o w   P o s i t i o n   c o m m a n d . 
 
 X 
 T h e   p o s i t i o n   o f   t h e   i t e m   o n   t h e   X   a x i s . 
 
 Y 
 T h e   p o s i t i o n   o f   t h e   i t e m   o n   t h e   Y   a x i s . 
 
 D X 
 T h e   c h a n g e   i n   X   a s   y o u   d r a w   o r   m o v e   a n   i t e m . 
 
 D Y 
 T h e   c h a n g e   i n   Y   a s   y o u   d r a w   o r   m o v e   a n   i t e m . 
 
 L e n 
 T h e   d i s t a n c e   b e t w e e n   t h e   s t a r t i n g   p o i n t   o f   t h e   o p e r a t i o n   a n d   t h e   c u r r e n t   p o s i t i o n . 
 
 A n g 
 T h e   a r c ,   i n   d e g r e e s ,   d e s c r i b e d   f r o m   t h e   s t a r t i n g   p o i n t   a s   y o u   d r a w   o r   m o v e   a n   i t e m . 
 
 
 P r e v i e w 
 D i s p l a y s   t h e   e n t i r e   i m a g e   i n   a   s e p a r a t e   P r e v i e w   W i n d o w . 
 
 I f   y o u   u s e   t h e   H a n d   T o o l   t o   p a n   t h r o u g h   a n   o v e r s i z e   i m a g e   i n   t h e   I m a g e   E d i t i n g   A r e a ,   t h e   a r e a   c u r r e n t l y   i n   t h e   I m a g e   E d i t i n g   A r e a   i s   o u t l i n e d   i n   t h e   P r e v i e w   W i n d o w . 
 
 Z o o m   I n 
 Z o o m   O u t 
 U s e   t h e s e   o p t i o n s   t o   m a g n i f y   o r   d e c r e a s e   t h e   m a g n i f i c a t i o n   o f   t h e   i m a g e   i n   t h e   I m a g e   E d i t i n g   A r e a . 
 
 
� F i l l   T o o l 
 
 U s e   t h e   F i l l   T o o l   t o   f i l l   a n y   e n c l o s e d   a r e a   o f   a n   i m a g e   w i t h   t h e   f o r e g r o u n d   c o l o r . 
 
 C l i c k   a n   e n c l o s e d   a r e a   o f   t h e   i m a g e   w i t h   t h e   F i l l   T o o l   t o   f i l l   t h e   a r e a   w i t h   t h e   f o r e g r o u n d   c o l o r .   
y� %����� |  &� " � � ����}� '���� ��
  ��  
[�   �= O p t i o n s   M e n u 
 
 T h e   O p t i o n s   M e n u   c o n t a i n s   t h e   f o l l o w i n g   o p t i o n s : 
 
 C h o o s e   F o n t . . . 
 O p e n s   a   f o n t   c h o o s e r . 
 
 U s e   t h e   f o n t   c h o o s e r   t o   s p e c i f y   f o n t   i n f o r m a t i o n   f o r   t e x t   a d d e d   t o   a n   i m a g e   w i t h   t h e   T e x t   T o o l . 
 
 E d i t   C o l o r s . . . 
 O p e n s   t h e   C o l o r   P a l e t t e   E d i t o r . 
 
 U s e   t h e   C o l o r   P a l e t t e   E d i t o r   t o   e d i t   t h e   c o l o r s   m a p p e d   t o   a n   i m a g e . 
 
 C r e a t e   T r a n s p a r e n c y 
 D e l e t e   T r a n s p a r e n c y 
 C r e a t e   T r a n s p a r e n c y   c r e a t e s   a   T r a n s p a r e n c y   E d i t i n g   A r e a .   D e l e t e   T r a n s p a r e n c y   r e m o v e s   a   p r e v i o u s l y   c r e a t e d   T r a n s p a r e n c y   E d i t i n g   A r e a . 
 
 I n   a   T r a n s p a r e n c y   E d i t i n g   A r e a   y o u   c r e a t e   a   t r a n s p a r e n c y ,   o r   m a s k ,   f o r   a n   i m a g e .   T r a n s p a r e n c i e s   a r e   u s e f u l   w h e n   f o r   i m a g e s   t h a t   n e e d s   t o   b e   v i s i b l e   a g a i n s t   v a r i o u s   b a c k g r o u n d s . 
 
 
[ D r o p p e r 
 
 U s e   t h e   D r o p p e r   T o o l   t o   p i c k   u p   t h e   c o l o r   f r o m   a   p i x e l . 
 
 C l i c k   a n y w h e r e   i n   t h e   I m a g e   E d i t i n g   A r e a   o r   t h e   C o l o r   P a l e t t e   t o   p i c k   u p   a   c o l o r .   T h e   c o l o r   y o u   p i c k   u p   i s   d i s p l a y e d   i n   t h e   F o r e g r o u n d   C o l o r   B o x . 
 
 T o   p i c k   u p   a   b a c k g r o u n d   c o l o r ,   p r e s s   t h e   C o n t r o l   k e y   w h e n   y o u   c l i c k   t h e   D r o p p e r   T o o l .   
����   �  �    (� P a l e E d S e t t i n g C o l o r s
[�   �
c�    9(� T o o l   P a l e t t e 
 
 T h e   T o o l   P a l e t t e   c o n t a i n s   t h e   f o l l o w i n g   i m a g e   e d i t i n g   t o o l s   f o r   d r a w i n g   i n   t h e   I m a g e   E d i t i n g   A r e a .   T h e   k e y b o a r d   m a c r o   f o r   e a c h   t o o l   i s   a l s o   l i s t e d . 
 
 
 H a n d   < H > 	 	 D r o p p e r   < D > 
 S e l e c t i o n   < S > 	 	 L a s s o   < S h i f t - S > 
 F i l l   < F > 	 	 S p r a y   C a n   T o o l   < A > 
 E r a s e r   < E > 	 	 T e x t   < T > 
 P e n c i l   < P > 	 	 L i n e   < L > 
 E l l i p s e   < E > 	 	 S o l i d   E l l i p s e   < S h i f t - C > 
 R e c t a n g l e < R > 	 	 S o l i d   R e c t a n g l e   < S h i f t - R > 
 
 
 T o   u s e   a   t o o l   f r o m   t h e   T o o l   P a l e t t e : 
 
 1 .   C l i c k   t h e   t o o l   y o u   w a n t   t o   u s e . 
 
 T h e   p o i n t e r   c h a n g e s   t o   t h e   a p p r o p r i a t e   c u r s o r   f o r   t h e   t o o l   y o u   s e l e c t e d .   
 
 2 .   C l i c k   a n d / o r   d r a g   t h e   p o i n t e r   i n   t h e   I m a g e   E d i t i n g   A r e a . 
 
 Y o u   c a n   a l s o   u s e   k e y b o a r d   m a c r o s   t o   s e l e c t   t o o l s   f r o m   t h e   T o o l   P a l e t t e . 
 
' S e l e c t i o n   T o o l 
 
 U s e   t h e   S e l e c t i o n   T o o l   t o   s e l e c t   a   r e c t a n g u l a r   a r e a   o f   a n   i m a g e   f o r   e d i t i n g . 
 
 D r a g   t h e   p o i n t e r   w i t h   t h e   S e l e c t i o n   T o o l   t o   d e s c r i b e   t h e   s e l e c t e d   a r e a   o f   t h e   i m a g e .   T o   s e l e c t   t h e   e n t i r e   I m a g e   E d i t i n g   A r e a ,   d o u b l e - c l i c k   t h e   S e l e c t i o n   T o o l   i n   t h e   T o o l   P a l e t t e .   
"a�����    x x##������NN4444==33"a            �  �    ) T o o l P a l e t t e ��
jz    �   //    �`   *   �( = K e y b o a r d   M a c r o s 
 
 K e y b o a r d   m a c r o s   p r o v i d e   a   s h o r t - c u t   f o r   s e l e c t i n g   t o o l s   f r o m   t h e   T o o l   P a l e t t e .   T h e y   a r e   u s e f u l   i f   y o u   w a n t   t o   s e l e c t   a   n e w   t o o l   w i t h o u t   l o s i n g   t h e   p o s i t i o n   o f   t h e   p o i n t e r   i n   t h e   I m a g e   E d i t i n g   A r e a . 
 
 K e y b o a r d   m a c r o s   f o r   i m a g e   e d i t i n g   t o o l s   a r e   c a s e - i n s e n s i t i v e . 
 
 T o   u s e   a   k e y b o a r d   m a c r o : 
 
 1 .   S e l e c t   t h e   I m a g e   E d i t i n g   A r e a   t o   g i v e   i t   f o c u s . 
 
 2 .   P r e s s   t h e   k e y   ( o r   k e y   c o m b i n a t i o n )   f o r   t h e   k e y b o a r d   m a c r o   y o u   w a n t . 
 
 T h e   c u r s o r   c h a n g e s   t o   r e f l e c t   t h e   n e w   e d i t i n g   t o o l . 
 
 N O T E :   F o r   o n e   t i m e   u s e   o f   a n   e d i t i n g   t o o l   u s e   t h e   A l t   k e y   m o d i f i e r   w i t h   t h e   k e y b o a r d   m a c r o .   A f t e r   d r a w i n g   w i t h   a   t o o l   s e l e c t e d   f o r   o n e   t i m e   u s e ,   t h e   c u r s o r   r e v e r t s   t o   t h e   p r e v i o u s   t o o l . 
 
; S p r a y   C a n   T o o l 
 
 U s e   t h e   S p r a y   C a n   T o o l   t o   d r a w   t h e   f o r e g r o u n d   c o l o r   w i t h   a   " s p r a y "   p a t t e r n . 
 
 D r a g   t h e   S p r a y   C a n   T o o l   a c r o s s   t h e   i m a g e   t o   d r a w   t h e   p a t t e r n .   
 T o o l P a l e t t eL  F  N V ] c k x { � � � � � � � � � � � � � � � � � � � �&-4
k5    	  
  �    + C o l o r P a l e t t e  C o l o r P a l P a l M e n u E d i t C o l o r P a l
kV   7  I n s t a l l C o l o r P a l
k|   v" C o l o r P a l F i l e M e n u
k� 	  �" C o l o r P a l E d i t M e n u�/� E r a s e r   T o o l 
 
 U s e   t h e   E r a s e r   T o o l   t o   r e p l a c e   t h e   c o l o r   o f   a n   i m a g e   w i t h   t h e   b a c k g r o u n d   c o l o r . 
 
 D r a g   t h e   E r a s e r   T o o l   o v e r   t h e   a r e a   y o u   w a n t   t o   e r a s e .   P r e s s   t h e   S h i f t   k e y   b e f o r e   e r a s i n g   t o   c o n s t r a i n   t h e   E r a s e r   T o o l   h o r i z o n t a l l y   o r   v e r t i c a l l y .   T o   c l e a r   t h e   e n t i r e   e d i t i n g   a r e a ,   c l i c k   i n   t h e   I m a g e   E d i t i n g   A r e a ,   a n d   t h e n   d o u b l e - c l i c k   t h e   E r a s e r   T o o l   i n   t h e   T o o l   P a l e t t e .   

k� 	  �  C o l o r P a l P a l M e n u
n�     C o l o r P a l B u t t o n s
o   
  �H   -   d�    �    ,%   C o l o r P a l P a l M e n u
oz      ] a) *('  ";;   �.P     � T e x t   T o o l 
 
 U s e   t h e   T e x t   T o o l   t o   p l a c e   t e x t   i n t o   t h e   i m a g e . 
 
 C l i c k   i n   t h e   I m a g e   E d i t i n g   A r e a   w i t h   t h e   T e x t   T o o l   t o   o p e n   a n   I m a g e   T e x t   W i n d o w .   T e x t   e n t e r e d   i n   t h e   I m a g e   T e x t   W i n d o w   a p p e a r s   a s   a   s e l e c t i o n   i n   t h e   i m a g e .   
� L i n e   T o o l 
 
 U s e   t h e   L i n e   T o o l   t o   d r a w   s t r a i g h t   l i n e s . 
 
 D r a g   t h e   L i n e   T o o l   i n   t h e   I m a g e   E d i t i n g   A r e a   t o   d r a w   a   s t r a i g h t   l i n e .   P r e s s   t h e   S h i f t   k e y   d u r i n g   t h e   d r a g   o p e r a t i o n   t o   c o n s t r a i n   t h e   l i n e   h o r i z o n t a l l y ,   v e r t i c a l l y ,   o r   t o   a   4 5 - d e g r e e   a n g l e .   

s� 	  "" #!   $  �    ." C o l o r P a l F i l e M e n u0,  0 O P e n c i l 
 
 U s e   t h e   P e n c i l   T o o l   t o   d r a w   o r   e r a s e   o n e   p i x e l   a t   a   t i m e . 
 
 C l i c k   i n   t h e   I m a g e   E d i t i n g   A r e a   w i t h   t h e   P e n c i l   T o o l   t o   d r a w   o r   e r a s e   a   p i x e l .   I f   t h e   P e n c i l   T o o l   i s   u s e d   o n   a n   i m a g e   a r e a   t h a t   c o n t a i n s   t h e   f o r e g r o u n d   c o l o r ,   t h e   P e n c i l   T o o l   d r a w s   t h e   b a c k g r o u n d   c o l o r .   O t h e r w i s e ,   t h e   P e n c i l   T o o l   d r a w s   t h e   f o r e g r o u n d   c o l o r . 
 
 D r a g   t h e   P e n c i l   T o o l   t o   d r a w   a   c o n t i n u o u s   l i n e .   U s e   F a t   B i t s   m o d e   t o   d r a w   o n e   p i x e l   a t   a   t i m e .   
   �?�kBp��  +  �    /
w�    @ E d i t C o l o r P a l3
{�   �"b"    � � � �[[	AAYY--	       2  �    0  � E l l i p s e   T o o l 
 
 U s e   t h e   E l l i p s e   T o o l   t o   d r a w   a n   e l l i p s e . 
 
 D r a g   t h e   E l l i p s e   T o o l   i n   t h e   I m a g e   E d i t i n g   A r e a   t o   d r a w   a n   e l l i p s e .   P r e s s   t h e   S h i f t   k e y   d u r i n g   t h e   d r a g   o p e r a t i o n   t o   c o n s t r a i n   t h e   e l l i p s e   t o   a   c i r c l e .   
� S o l i d   E l l i p s e   T o o l 
 
 U s e   t h e   S o l i d   E l l i p s e   T o o l   t o   d r a w   a   s o l i d   e l l i p s e . 
 
 D r a g   t h e   S o l i d   E l l i p s e   T o o l   i n   t h e   I m a g e   E d i t i n g   A r e a   t o   d r a w   a   s o l i d   e l l i p s e .   P r e s s   t h e   S h i f t   k e y   d u r i n g   t h e   d r a g   o p e r a t i o n   t o   c o n s t r a i n   t h e   e l l i p s e   t o   a   c i r c l e .   
0 1/.((**  C o l o r P a l B u t t o n s
  �    1  **99�7 865!e1  �� �� �       � R e c t a n g l e   T o o l 
 
 U s e   t h e   R e c t a n g l e   T o o l   t o   d r a w   a   r e c t a n g l e . 
 
 D r a g   t h e   R e c t a n g l e   T o o l   i n   t h e   I m a g e   E d i t i n g   A r e a   t o   d r a w   a   r e c t a n g l e .   P r e s s   t h e   S h i f t   k e y   d u r i n g   t h e   d r a g   o p e r a t i o n   t o   c o n s t r a i n   t h e   r e c t a n g l e   t o   a   s q u a r e .   
� S o l i d   R e c t a n g l e   T o o l 
 U s e   t h e   S o l i d   R e c t a n g l e   T o o l   t o   d r a w   a   s o l i d   r e c t a n g l e . 
 
 D r a g   t h e   S o l i d   R e c t a n g l e   T o o l   i n   t h e   I m a g e   E d i t i n g   A r e a   t o   d r a w   a   s o l i d   r e c t a n g l e .   P r e s s   t h e   S h i f t   k e y   d u r i n g   t h e   d r a g   o p e r a t i o n   t o   c o n s t r a i n   t h e   r e c t a n g l e   t o   a   s q u a r e .   
Q                                                                                � C o l o r   P a l e t t e 
 
 T h e   C o l o r   P a l e t t e   c o n t a i n s   1 6   c o l o r s   r e a d i l y   a v a i l a b l e   t o   u s e   i n   y o u r   i m a g e .   T h e   1 6   c o l o r s   o n   t h e   C o l o r   P a l e t t e   r e p r e s e n t   t h e   m o s t   r e c e n t l y   u s e d   c o l o r s   f r o m   t h e   E x t e n d e d   C o l o r   P a l e t t e . 
 
 T h e   C o l o r   P a l e t t e   i s   l o c a t e d   b e t w e e n   t h e   T o o l   P a l e t t e   a n d   t h e   I m a g e   E d i t i n g   A r e a . 
 
 E x t e n d e d   C o l o r   P a l e t t e 
 
 T h e   E x t e n d e d   C o l o r   P a l e t t e   r e p r e s e n t s   t h e   c o m p l e t e   c o l o r   p a l e t t e   i n s t a l l e d   w i t h   t h e   i m a g e .   T h i s   p a l e t t e   c o n t a i n s   u p   t o   2 5 6   c o l o r s .   U s e   t h e   C o l o r   P a l e t t e   E d i t o r   t o   e d i t   c o l o r s   o n   t h e   E x t e n d e d   C o l o r   P a l e t t e   o r   t o   i n s t a l l   d i f f e r e n t   c o l o r   p a l e t t e s . 
 
 T o   v i e w   t h e   E x t e n d e d   C o l o r   P a l e t t e ,   c l i c k   a n d   h o l d   o n   e i t h e r   t h e   F o r e g r o u n d   o r   B a c k g r o u n d   C o l o r   B o x . 
 
 F o r e g r o u n d   C o l o r   B o x 
 B a c k g r o u n d   C o l o r   B o x 
 
 B e n e a t h   t h e   C o l o r   P a l e t t e   a r e   t h e   F o r e g r o u n d   C o l o r   B o x   a n d   t h e   B a c k g r o u n d   C o l o r   B o x .   ( T h e   F o r e g r o u n d   C o l o r   B o x   i s   t o   t h e   r i g h t   a n d   i n   f r o n t   o f   t h e   B a c k g r o u n d   C o l o r   B o x . ) 
 
 U s e   t h e   C o l o r   P a l e t t e ,   F o r e g r o u n d   C o l o r   B o x ,   a n d   B a c k g r o u n d   C o l o r   b o x   t o   s e t   c o l o r s   f o r   d r a w i n g . 
 
 
i                                                                                                        _ S e t t i n g   C o l o r s   f o r   D r a w i n g 
 
 T h e   f o l l o w i n g   t o o l s   f r o m   t h e   T o o l   P a l e t t e   u s e   f o r e g r o u n d   a n d   b a c k g r o u n d   c o l o r s   f o r   d r a w i n g : 
 
 * 	 S p r a y   C a n   T o o l 
 * 	 P e n c i l   T o o l 
 * 	 L i n e   T o o l 
 * 	 E l l i p s e   T o o l s 
 * 	 R e c t a n g l e   T o o l s 
 
 
 U s e   a n y   o f   t h e   f o l l o w i n g   m e t h o d s   t o   s e t   t h e   f o r e g r o u n d   a n d   b a c k g r o u n d   c o l o r s   f o r   d r a w i n g . 
 
 T o   s e t   t h e   f o r e g r o u n d   c o l o r   u s i n g   t h e   C o l o r   P a l e t t e : 
 
 1 .   C l i c k   o n   a   c o l o r   i n   t h e   C o l o r   P a l e t t e . 
 
 T h e   c o l o r   i s   d i s p l a y e d   i n   t h e   F o r e g r o u n d   C o l o r   B o x .   C o l o r s   c a n   b e   s e t   b e f o r e   o r   a f t e r   c l i c k i n g   o n   a   d r a w i n g   t o o l . 
 
 
 T o   s e t   t h e   b a c k g r o u n d   c o l o r   u s i n g   t h e   C o l o r   P a l e t t e : 
 
 1 .   P r e s s   t h e   C o n t r o l   k e y   a n d   c l i c k   o n   a   c o l o r   i n   t h e   C o l o r   P a l e t t e .   
 
 T h e   c o l o r   i s   d i s p l a y e d   i n   t h e   B a c k g r o u n d   C o l o r   B o x .   C o l o r s   c a n   b e   s e t   b e f o r e   o r   a f t e r   c l i c k i n g   o n   a   d r a w i n g   t o o l . 
 
 
 T o   s e t   t h e   f o r e g r o u n d   c o l o r   u s i n g   t h e   E x t e n d e d   C o l o r   P a l e t t e : 
 
 1 .   C l i c k   a n d   h o l d   t h e   F o r e g r o u n d   C o l o r   B o x . 
 
 T h e   e x t e n d e d   C o l o r   P a l e t t e   i s   d i s p l a y e d .   T h e   c u r r e n t   f o r e g r o u n d   c o l o r   i s   i n d i c a t e d   i n   t h e   p a l e t t e . 
 
 2 .   D r a g   t h e   p o i n t e r   t o   a   c o l o r   i n   t h e   E x t e n d e d   C o l o r   P a l e t t e   a n d   r e l e a s e   t h e   p o i n t e r . 
 
 T h e   f o r e g r o u n d   c o l o r   i s   s e t   t o   t h e   c o l o r   y o u   s e l e c t e d .   T h e   c o l o r   i s   d i s p l a y e d   i n   t h e   F o r e g r o u n d   C o l o r   B o x   a n d   i s   a d d e d   t o   t h e   C o l o r   P a l e t t e . 
 
 S i m i l a r l y ,   t h e   b a c k g r o u n d   c o l o r   c a n   b e   s e t   f r o m   t h e   B a c k g r o u n d   C o l o r   B o x . 
 
 
 T o   s e t   t h e   f o r e g r o u n d   c o l o r   u s i n g   t h e   D r o p p e r   T o o l : 
 
 1 .   S e l e c t   t h e   D r o p p e r   T o o l   f r o m   t h e   T o o l   P a l e t t e . 
 
 T h e   c u r s o r   c h a n g e s   t o   a n   e y e - d r o p p e r . 
 
 2 .   W i t h   t h e   D r o p p e r   T o o l ,   s e l e c t   a   c o l o r   i n   t h e   I m a g e   E d i t i n g   A r e a ,   o r   f r o m   t h e   C o l o r   P a l e t t e . 
 
 T h e   f o r e g r o u n d   c o l o r   i s   s e t   t o   t h e   c o l o r   o f   t h e   p i x e l   y o u   s e l e c t e d   a n d   i s   d i s p l a y e d   i n   t h e   F o r e g r o u n d   C o l o r   B o x . 
 
 T o   s e t   t h e   b a c k g r o u n d   c o l o r ,   p r e s s   t h e   C o n t r o l   k e y   w h i l e   s e l e c t i n g   a   c o l o r   w i t h   t h e   D r o p p e r   T o o l . 
 
 
_ L i n e   W i d t h   P a l e t t e 
 
 U s e   t h e   L i n e   W i d t h   P a l e t t e   t o   s e t   t h e   l i n e   w i d t h   f o r   d r a w i n g .   S e t t i n g   t h e   l i n e   w i d t h   a p p l i e s   t o   t h e   f o l l o w i n g   d r a w i n g   t o o l s   f r o m   t h e   T o o l   P a l e t t e : 
 
 * 	 L i n e   T o o l 
 * 	 E l l i p s e   T o o l s 
 * 	 R e c t a n g l e   T o o l s 
 
 
 
 T o   s e t   t h e   l i n e   w i d t h ,   u s e   t h e   p o i n t e r   t o   s e l e c t   o n e   o f   t h e   f o u r   w i d t h s   a v a i l a b l e . 
 
 
?                                                              G C o l o r   P a l e t t e   E d i t o r 
 
 E a c h   i m a g e   i n   t h e   I m a g e   E d i t o r   h a s   a n   a s s o c i a t e d   c o l o r   p a l e t t e   c o n t a i n i n g   u p   t o   2 5 6   c o l o r s .   T h i s   c o l o r   p a l e t t e   i s   t h e   " E x t e n d e d   C o l o r   P a l e t t e "   y o u   c a n   v i e w   f r o m   e i t h e r   t h e   F o r e g r o u n d   o r   B a c k g r o u n d   C o l o r   B o x   i n   t h e   I m a g e   E d i t o r . 
 
 U s e   t h e   C o l o r   P a l e t t e   E d i t o r   t o   l o a d   a   n e w   c o l o r   p a l e t t e   o r   e d i t   a   c o l o r   p a l e t t e .   A f t e r   l o a d i n g   o r   e d i t i n g   a   c o l o r   p a l e t t e   i n s t a l l   t h e   n e w   c o l o r   p a l e t t e   t o   a p p l y   i t   t o   t h e   c u r r e n t   i m a g e . 
 
 T h e   C o l o r   P a l e t t e   E d i t o r   h a s   t h e   f o l l o w i n g   c o m p o n e n t s : 
 
 F i l e   M e n u 
 E d i t   M e n u 
 P a l e t t e s   M e n u 
 E d i t i n g   B u t t o n s 
 
# C o l o r   P a l e t t e   E d i t o r   E d i t   M e n u 
 
 T h e   C o l o r   P a l e t t e   E d i t   M e n u   c o n t a i n s   t h e   f o l l o w i n g   o p t i o n s : 
 
 U n d o   S e t   I m a g e 
 T h e   U n d o   S e t   I m a g e   o p t i o n   u n i n s t a l l s   p r e v i o u s l y   i n s t a l l e d   c o l o r   p a l e t t e s .   T h i s   o p t i o n   o n l y   u n i n s t a l l s   i m a g e s   t h a t   h a v e   b e e n   i n s t a l l e d   d u r i n g   t h e   c u r r e n t   e d i t i n g   s e s s i o n . 
 
 C u t 
 C o p y 
 P a s t e 
 U s e   t h e s e   o p t i o n s   t o   p e r f o r m   e d i t i n g   a c t i o n s   o n   c o l o r s   s e l e c t e d   f o r   e d i t i n g   i n   t h e   C o l o r   P a l e t t e   E d i t o r . 
 
 �                                                                                                                                                 � C o l o r   P a l e t t e   E d i t o r   F i l e   M e n u 
 
 T h e   C o l o r   P a l e t t e   E d i t o r   F i l e   M e n u   c o n t a i n s   t h e   f o l l o w i n g   o p t i o n s : 
 
 R e v e r t 
 R e s t o r e s   t h e   C o l o r   P a l e t t e   E d i t o r   t o   t h e   l a s t   i n s t a l l e d   v e r s i o n .   A l l   c h a n g e s   m a d e   t o   t h e   e d i t o r   s i n c e   t h e   l a s t   v e r s i o n   a r e   l o s t . 
 
 N o t e   t h a t   s a v i n g   a   c o l o r   p a l e t t e   d o e s   n o t   i n s t a l l   t h e   p a l e t t e .   Y o u   c a n   s t i l l   r e v e r t   t h e   C o l o r   P a l e t t e   E d i t o r   t o   t h e   i n s t a l l e d   v e r s i o n   a f t e r   s a v i n g   a   c o l o r   p a l e t t e . 
 
 S a v e . . . 
 S a v e s   t h e   c o l o r   p a l e t t e   c u r r e n t l y   b e i n g   e d i t e d . 
 
 S a v e d   p a l e t t e s   a r e   a v a i l a b l e   a c r o s s   d i f f e r e n t   e d i t i n g   s e s s i o n s .   U s e   t h e   P a l e t t e s   M e n u   t o   l o a d   s a v e d   p a l e t t e s   i n t o   t h e   C o l o r   P a l e t t e   E d i t o r .   
 
 � /
	
# &#(,E. � 	AttributeContextqBlock!untQsExtraKeywordBlockLengthasinkListAType	NodeBlockADataA	TextsOffsetasTagextAAttributes	itleQs
ypeVersionvhelpDocument �    >   � 6    �  �   � >  >      �   ` H  � � �   �      	Sk  A � �5 K � �                                                                                                                                                                                           � C o l o r   P a l e t t e   E d i t o r   P a l e t t e s   M e n u 
 
 U s e   t h e   P a l e t t e s   M e n u   t o   l o a d   c o l o r   p a l e t t e s   i n t o   t h e   C o l o r   P a l e t t e   E d i t o r . 
 
 T h e   f o l l o w i n g   o p t i o n s   a r e   a v a i l a b l e   f r o m   t h e   P a l e t t e s   M e n u : 
 
 D e l e t e 
 D e l e t e   a   p r e v i o u s l y   s a v e d   p a l e t t e . 
 
 P a l e t t e s   a r e   s a v e d   w i t h   t h e   S a v e . . .   o p t i o n   f r o m   t h e   C o l o r   P a l e t t e   E d i t o r   F i l e   M e n u . 
 
 D e f a u l t   P a l e t t e   L i s t 
 T h i s   i s   a   l i s t   o f   c o l o r   p a l e t t e s   t h a t   a r e   a l w a y s   a v a i l a b l e   f r o m   t h e   C o l o r   P a l e t t e   E d i t o r .   S e l e c t   a   p a l e t t e   f r o m   t h i s   l i s t   t o   l o a d   t h e   p a l e t t e   i n t o   t h e   C o l o r   P a l e t t e   E d i t o r . 
 
 T h e   c o l o r   p a l e t t e s   a v a i l a b l e   a r e : 
 
 * 	 E G A   P a l e t t e 
 * 	 E a r t h   T o n e s 
 * 	 H u e s   1 6 
 * 	 P a s t e l s 
 * 	 R a i n b o w 
 
 
 S a v e d   P a l e t t e   L i s t 
 T h i s   i s   a   l i s t   o f   p r e v i o u s l y   s a v e d   p a l e t t e s .   S e l e c t   a   p a l e t t e   f r o m   t h i s   l i s t   t o   l o a d   t h e   p a l e t t e   i n t o   t h e   C o l o r   P a l e t t e   E d i t o r . 
 
3                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 � C o l o r   P a l e t t e   E d i t i n g   B u t t o n s 
 
 U s e   t h e   C o l o r   P a l e t t e   B u t t o n s   t o   e d i t   c o l o r s   o n   t h e   p a l e t t e . 
 
 T h e   f o l l o w i n g   b u t t o n s   a r e   a v a i l a b l e   t o   e d i t   a   c o l o r   ( o r   s e r i e s   o f   c o l o r s ) : 
 
 N e w 
 A d d s   a   n e w   c o l o r   t o   t h e   p a l e t t e .   Y o u   c a n   k e e p   a d d i n g   c o l o r s   u n t i l   t h e   p a l e t t e   c o n t a i n s   2 5 6   c o l o r s . 
 
 D e l e t e 
 R e m o v e s   t h e   s e l e c t e d   c o l o r   o r   c o l o r s . 
 
 P i c k . . . 
 O p e n s   a   c o l o r   c h o o s e r .   R e d e f i n e   t h e   s e l e c t e d   c o l o r   w i t h   t h e   c o l o r   c h o o s e r . 
 
 N o t e   t h a t   d o u b l e - c l i c k i n g   o n   a   c o l o r   a l s o   o p e n s   t h e   c o l o r   c h o o s e r   t o   e d i t   t h e   c o l o r . 
 
 R a m p 
 C r e a t e s   a   r a n g e   o f   c o l o r s   f r o m   w h i t e   t o   b l a c k .   T h e   f i r s t   c o l o r   i n   t h e   o r i g i n a l   s e r i e s   b e c o m e s   t h e   m i d d l e   c o l o r   o f   t h e   r a m p . 
 
 B l e n d 
 M o d i f i e s   a   s e r i e s   o f   c o l o r s   s o   t h a t   t h e   c o l o r s   r a n g e   g r a d u a l l y   f r o m   t h e   f i r s t   c o l o r   i n   t h e   o r i g i n a l   s e r i e s   t o   t h e   l a s t   c o l o r   i n   t h e   o r i g i n a l   s e r i e s . 
 
 C o n t r a s t 
 C h a n g e s   t h e   s e l e c t e d   c o l o r ( s )   t o   i t s   c o m p l e m e n t . 
 
 L i g h t e r 
 A d d s   w h i t e   t o   t h e   s e l e c t e d   c o l o r ( s ) . 
 
 D a r k e r 
 A d d s   b l a c k   t o   t h e   s e l e c t e d   c o l o r ( s ) . 
 
 W a r m e r 
 A d d s   r e d   t o   t h e   s e l e c t e d   c o l o r ( s ) . 
 
 C o o l e r 
 A d d s   b l u e   t o   t h e   s e l e c t e d   c o l o r ( s ) . 
 
                  � E d i t i n g   a   C o l o r   P a l e t t e 
 
 I n   t h e   C o l o r   P a l e t t e   E d i t o r ,   b e f o r e   y o u   c a n   e d i t   a   c o l o r   o n   a   c o l o r   p a l e t t e ,   y o u   m u s t   f i r s t   s e l e c t   t h e   c o l o r . 
 
 T o   s e l e c t   a   c o l o r   o r   s e r i e s   o f   c o l o r s   d o   e i t h e r   o f   t h e   f o l l o w i n g : 
 
 * 	 C l i c k   o n   t h e   c o l o r   i n   t h e   c o l o r   p a l e t t e . 
 
 * 	 D r a g   t h e   p o i n t e r   o v e r   a   s e r i e s   o f   c o l o r s . 
 
 S e l e c t e d   c o l o r s   a p p e a r   o u t l i n e d   i n   t h e   c o l o r   p a l e t t e . 
 
 T o   e d i t   s e l e c t e d   c o l o r s   o n   t h e   c o l o r   p a l e t t e : 
 
 1 .   C l i c k   o n   o n e   o f   t h e   e d i t i n g   b u t t o n s . 
 
 T h e   e d i t i n g   b u t t o n s   p r o v i d e   v a r i o u s   o p t i o n s   f o r   e d i t i n g   c o l o r s . 
 
                  	� I n s t a l l i n g   a   C o l o r   P a l e t t e 
 
 A f t e r   l o a d i n g   o r   e d i t i n g   a   c o l o r   p a l e t t e   i n   t h e   C o l o r   P a l e t t e   E d i t o r ,   y o u   n e e d   t o   i n s t a l l   t h e   c o l o r   p a l e t t e . 
 
 I n s t a l l i n g   t h e   c o l o r   p a l e t t e   m a p s   t h e   p a l e t t e   t o   t h e   i m a g e   c u r r e n t l y   b e i n g   e d i t e d   i n   t h e   I m a g e   E d i t o r .   I t   a l s o   m a k e s   t h e   c o l o r   p a l e t t e   a v a i l a b l e   f o r   d r a w i n g . 
 
 
 T o   i n s t a l l   a   c o l o r   p a l e t t e   f o r   a n   i m a g e : 
 
 1 .   A f t e r   l o a d i n g   o r   e d i t i n g   a   c o l o r   p a l e t t e ,   c l i c k   o n   t h e   I n s t a l l   B u t t o n . 
 
 T h e   c o l o r   p a l e t t e   i s   i n s t a l l e d .   T h e   C o l o r   P a l e t t e   E d i t o r   c l o s e s   a n d   t h e   i m a g e   i n   t h e   I m a g e   E d i t o r   c h a n g e s   t o   r e f l e c t   t h e   n e w l y   i n s t a l l e d   c o l o r   p a l e t t e . 
 
 
 T o   u n i n s t a l l   a   c o l o r   p a l e t t e   f o r   a n   i m a g e : 
 
 1 .   F r o m   t h e   E d i t   M e n u ,   s e l e c t   U n d o   S e t   I m a g e . 
 
 T h e   i m a g e   i n   t h e   I m a g e   E d i t o r   i s   s e t   t o   t h e   p r e v i o u s l y   i n s t a l l e d   c o l o r   p a l e t t e . 
 
 
 R e m a p   T o   C l o s e s t   C o l o r 
 W h e n   c o l o r   p a l e t t e s   a r e   i n s t a l l e d   f o r   a n   i m a g e ,   t h e   c o l o r s   o f   t h e   n e w l y   i n s t a l l e d   p a l e t t e   a r e   m a t c h e d   t o   t h e   c l o s e s t   c o l o r s   o n   t h e   p r e v i o u s   i n s t a l l e d   c o l o r   p a l e t t e .   T h i s   d e f a u l t   b e h a v i o r   m i n i m i z e s   c h a n g e s   t o   a n   i m a g e   w h e n   i n s t a l l i n g   a   n e w   p a l e t t e . 
 
 Y o u   c a n   o v e r r i d e   t h i s   d e f a u l t   b e h a v i o r   b y   u n s e l e c t i n g   t h e   R e m a p   t o   C l o s e s t   C o l o r   t o g g l e .   W h e n   R e m a p   T o   C l o s e s t   C o l o r   i s   n o t   s e l e c t e d ,   c o l o r s   o n   t h e   n e w l y   i n s t a l l e d   p a l e t t e   a r e   m a p p e d   a c c o r d i n g   t o   t h e i r   p o s i t i o n   o n   t h e   p a l e t t e . 
I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       
��8qr b
�ab�!B�ar �
ab�qb5Ab�q"caabhbarj�(a",(ab�&q"�&aNb\&aV"�&!]r�&!cB�&akrlaxb^&q{b+�&b �+�b& �"8�&r �:�b& �";&" �;r& �b;u&r �;�"& �b;�&" �;�b& �rCx& �C�b& �bC�&b �C�"& �bC�&b �S�r& �bS�&r �S�"& �r[�&r �cE"& �bc�&rj�r&rom&"o�b&"s�&r&o�b&-r{�&b4{�b&
�b2a2aZ"2#A2b�a"5,a7rh,!7"�,!7b�,a7"�,a7b
�,q7b�,a7b�,q7"�,a7b�,a7",a7bB,a7bd,a7b~,a7r�abG,7�a"�qrea"�ab`q"B,aLb�(a"d,qL"!bAabR2Ab�qN"",aTb�(a"�!b�qb�!btab:!Vrm,a[r�!"|,a[b�ab�ab�ar�aby(qr�a"�Qb�ab>q"�acb�,ah",!hbS(qb�,ahb1QbyAb�q"�abeak"�,aqr�,!qb�,qqb#�,aqb*M,qqb*w,aqb*�.a"�,!qr�,!B+s(ab#�ab+�q"+�ab+�q"/!{rt,b �/<r(/xb, �b/`q"/kqr+�ab�ab�r �+~b, �r/�," �/�(8�r, �b/�ab/�a"+�ab8�qb/�r �8�", �r9,b �9Bb, �b9^, �9~", �b9�,r �9�", �b9�,B �9�r, �r:,b �:,", �b:H,R �:j", �b:�," �:�R, �":�ab8�,b �9$r:�B/�b:�b:�":�r�r:�b:�r:�b(;'r:�r;b;b:�r �b;,r �;Z";QR;r;j";0r;e";nb;}b;�b;�r;�b;�b;�r;�b;�b;�";�";�b;�b;�b;�b;�r ;�" ;�" ;�b ;�b;�b!;�"!C�b!;�"!C�"C�b"C�""C�r"C�b"C�bC�b#C�r#C�b#C�b#C�bC�r$C�b$C�b$C�"$C�bSzb%C�r%S�R%S�"%C�bS�"&C�b&S�r&S�b&S�rS�b'S�b'S�r'S�b'S�b([�r(S�"(S�r(S�b(S�b �bS�,r �S�b(c�", �R[�!)bcN!)bcgq)rcua)"c~b �[�b, �b[�(q"c�a*bc�a*rc�q*"c@q*bc�b �[�b,rc�(!Rj�a+ra+"!a+rq+"bk",
b,b
kqR,
bk�,b
k�r,
bn�,b
ob,
"o:(aboY,b
j�b,oPr,c�b,%",S�brc�,bo�boEb-o�"-o�r-[�b-c�b(s�r.o�r.o�b.o�b.o�bboh,b$s�b(wwb/w^r/wPr/k�"/s�r&"s�,b+w�r(w�0w�0w�0w�0w�-bw�,2w��{�1{�b1{�1{��1s��