��       Td  b@b � F o n t   C h o o s e r"j" T h e   F o n t   C h o o s e r���,�� ��  ��   ��   ��   ��   ��   ����$ F o n t   D i s p l a y   A r e a* T y p e f a c e   F a m i l y   L i s t F a c e   L i s t2 S i z e   T e x t   F i e l d   a n d   L i s t P � � �S~* C o n f i r m a t i o n   B u t t o n s> S p e c i f y i n g   F o n t s   a n d   T y p e f a c e sG<    v f o n t c h s r��	 ;Na��� S i z e L i s t F a m i l y L i s t S p e c i f y F o n t s F a c e L i s t O v e r v i e w C o n f i r m B u t t o n s* I m a g e E d i t o r v f o n t c h s r( v s t y l e c h s r v f o n t c h s r D i s p l a y A r e a    *   f o n t   c h o o s e r	 "l�     S p e c i f y F o n t s��
K    & D i s p l a y A r e a
z   � F a m i l y L i s t
�   � F a c e L i s t
� 	  � S i z e L i s t
�   �!� F o n t   C h o o s e r 
 
 U s e   t h e   F o n t   C h o o s e r   t o   s p e c i f y   f o n t s   a n d   t y p e f a c e s   i n   y o u r   a p p l i c a t i o n . 
 
 T h e   F o n t   C h o o s e r   h a s   t h e   f o l l o w i n g   c o m p o n e n t s : 
 
 F o n t   D i s p l a y   A r e a 
 T y p e f a c e   F a m i l y   L i s t 
 F a c e   L i s t 
 S i z e   T e x t   F i e l d   a n d   L i s t 
 C o n f i r m a t i o n   B u t t o n s 
 
 C o n f i r m B u t t o n s
�   � � T h e   F o n t   D i s p l a y   A r e a   d i s p l a y s   a n   e x a m p l e   o f   t h e   c u r r e n t l y   s e l e c t e d   f o n t . 
 
 � T h e   T y p e f a c e   F a m i l y   L i s t   d i s p l a y s   t h e   t y p e f a c e s   a v a i l a b l e   o n   y o u r   s y s t e m . 
 
 � T h e   F a c e   L i s t   d i s p l a y s   t h e   f a c e s   a v a i l a b l e   f o r   t h e   f o n t   f a m i l y   s e l e c t e d   i n   t h e   F a m i l y   L i s t . 
 
2 	� � T h e   S i z e   L i s t   d i s p l a y s   t h e   s i z e s   a v a i l a b l e   f o r   t h e   c u r r e n t l y   s e l e c t e d   f o n t   f a m i l y . 
 
 U s e   t h e   S i z e   T e x t   F i e l d   t o   s p e c i f y   a   c u s t o m   s i z e   f o r   t h e   c u r r e n t   s e l e c t i o n .   W h e n   s i z e s   t h a t   a r e   n o t   i n   t h e   l i s t   a r e   s p e c i f i e d ,   t h e   n e w   s i z e   i s   a d d e d   t o   t h e   l i s t . 
 
~ U s e   t h e   c o n f i r m a t i o n   b u t t o n s   t o   a p p l y   t h e   c u r r e n t   s e l e c t i o n . 
 
  !	#"!#$"! � a-q!qaa
!aaaqaa	
aAaaa!qq!aqq!Aaa!a &qq(q,a� �"
�B �` ` qab �&� �                                                                                                                                        � T o   s p e c i f y   a   f o n t   a n d   t y p e f a c e : 
 
 1 .   S e l e c t   a   t y p e f a c e   f a m i l y ,   f a c e ,   a n d   s i z e   f r o m   t h e   l i s t s   i n   t h e   F o n t   C h o o s e r .   Y o u   c a n   a l s o   u s e   t h e   S i z e   t e x t   f i e l d   t o   s p e c i f y   a   s i z e . 
 
 Y o u r   s e l e c t i o n   i s   p r e v i e w e d   i n   t h e   F o n t   D i s p l a y   A r e a . 
 
 
 2 .   A p p l y   y o u r   s e l e c t i o n   w i t h   t h e   a p p r o p r i a t e   c o n f i r m a t i o n   b u t t o n s . 
 
 Y o u r   f o n t   s p e c i f i c a t i o n s   a r e   a p p l i e d   t o   y o u r   p r e v i o u s l y   s e l e c t e d   t e x t . 
 
 
 
 
 
 
 
 
 �q`aq�	AttributeAContextaqBlocka!untQsExtraKeywordBlockaLengthaasinkListATypeq	NodeBlockADataaA	TextsqOffsetAasqTagAextaAAttributesa	itleaQs
ypeVersionvhelpDocument$                                    1$p�b�"Bb}
aaE"ab�1xaasb&!r(ab9a"fab�!"�ab�ab�&qb
�&!b1a!"r&bJ!b!qbB,Abo,!B�,ar�,!"�,q"�a"*,qb�qbkab
var
{qb
q�