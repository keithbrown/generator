��     D  .�  6Ww   F i l e   C h o o s e r��� F i l e   C h o o s e rB b�� ��  ��      ����     ��  ����  ��   �� 	  �� 
  ��   ��   ��   ��   ��   ����6 N a v i g a t i n g   t h e   F i l e   S y s t e m H i s t o r y   M e n u" S �Y�����0Sh���. U s i n g   t h e   H i s t o r y   M e n u S p e c i a l   M e n u M a r k   P r o c e d u r e" U n m a r k   P r o c e d u r e V i e w   M e n u F i l t e r s   M e n u V o l u m e s   M e n u" P a t h   P o p - u p   M e n u F i l e   L i s t A r r o w   B u t t o n s* P a t h   N a m e   T e x t   F i e l d* C o n f i r m a t i o n   B u t t o n s4 R e s i z i n g   t h e   F i l e   C h o o s e r C o n f i r m B u t t o n s&bu����� >Wp�����o�p0)�E� O v e r v i e w R e s i z e U n m a r k P r o c P a t h M e n u F i l e L i s t* I m a g e E d i t o r v f i l e c h s r V i e w M e n u  v f i l e c h s r( H i s t o r y N a v i g a t e P r o c V o l u m e s M e n u H i s t o r y M e n u N a v i g a t e F i l e s F i l t e r s M e n u M a r k P r o c S p e c i a l M e n u A r r o w B u t t o n s P a t h F i e l d    *   f i l e   c h o o s e r.;EKSY^chmrw|�� ! "  #/$%&'()*+,-"b N a v i g a t e F i l e s2310 
i !   * H i s t o r y M e n u
�    � S p e c i a l M e n u
�    � V i e w M e n u
� 	   � F i l t e r s M e n u
     � V o l u m e s M e n u
$    � P a t h M e n u
H    � F i l e L i s t
f 	   � A r r o w B u t t o n s
�    � P a t h F i e l d
�    C o n f i r m B u t t o n s
�    R e s i z e
� /  ` jj  L L    4  	5<6789: H i s t o r y M e n u8 
F    � H i s t o r y M e n u
s    � P a t h M e n u
�   " A r r o w B u t t o n s
�   � F i l e L i s t
� 	  � ' T h e   F i l e   C h o o s e r 
 
 U s e   t h e   F i l e   C h o o s e r   t o   n a v i g a t e   t h r o u g h   y o u r   f i l e   s y s t e m   w h e n   o p e n i n g   o r   s a v i n g   f i l e s . 
 
 T h e   F i l e   C h o o s e r   h a s   t h e   f o l l o w i n g   c o m p o n e n t s : 
 
 H i s t o r y   M e n u 
 S p e c i a l   M e n u 
 V i e w   M e n u 
 F i l t e r s   M e n u 
 V o l u m e s   M e n u 
 P a t h   P o p - u p   M e n u 
 F i l e   L i s t 
 A r r o w   B u t t o n s 
 P a t h   N a m e   T e x t   F i e l d 
 C o n f i r m a t i o n   B u t t o n s 
 
 Y o u   c a n   r e s i z e   t h e   F i l e   C h o o s e r   ( m a k e   i t   w i d e r )   t o   d i s p l a y   m o r e   t h a n   o n e   d i r e c t o r y   l e v e l   a t   a   t i m e . 
 
 F i l e L i s t
( 	  � P a t h F i e l d
F   t   ��?@>= A  BFCD O( H i s t o r y N a v i g a t e P r o cH!	 
�   . M a r k P r o c
�  V
   f
+  � N a v i g a t i n g   t h e   F i l e   S y s t e m 
 
 T o   n a v i g a t e   y o u r   f i l e   s y s t e m   w i t h   t h e   F i l e   C h o o s e r ,   d o   o n e   o f   t h e   f o l l o w i n g : 
 
 * 	 S e l e c t   a   p a t h   f r o m   t h e   H i s t o r y   L i s t   i n   t h e   H i s t o r y   M e n u . 
 
 * 	 S e l e c t   a   p a t h   f r o m   t h e   M a r k e d   D i r e c t o r i e s   L i s t   i n   t h e   H i s t o r y   M e n u . 
 
 * 	 S e l e c t   a   c o m p o n e n t   f r o m   t h e   c u r r e n t   p a t h   u s i n g   t h e   P a t h   P o p - u p   M e n u . 
 
 * 	 M o v e   u p   o r   d o w n   a   l e v e l   f r o m   t h e   c u r r e n t l y   s p e c i f i e d   d i r e c t o r y   u s i n g   t h e   A r r o w   B u t t o n s . 
 
 * 	 D o u b l e - c l i c k   o n   a   d i r e c t o r y   o r   f i l e   i n   t h e   F i l e   L i s t . 
 
 * 	 S e l e c t   a   d i r e c t o r y   o r   f i l e   i n   t h e   F i l e   L i s t   a n d   a c c e p t   t h e   e n t r y   w i t h   t h e   p r o p e r   c o n f i r m a t i o n   b u t t o n   ( o r   p r e s s   E n t e r   t o   a c c e p t   t h e   e n t r y . ) 
 
 * 	 S p e c i f y   a   p a t h   n a m e   i n   t h e   P a t h   N a m e   F i e l d . 
 
 
 S p e c i a l M e n u U n m a r k P r o c� T o   c h a n g e   d i r e c t o r i e s   u s i n g   t h e   H i s t o r y   M e n u : 
 
 1 .   S e l e c t   a   n e w   d i r e c t o r y   f r o m   e i t h e r   t h e   H i s t o r y   L i s t   o r   t h e   M a r k e d   D i r e c t o r i e s   L i s t . 
 
 T h e   d i r e c t o r y   d i s p l a y e d   i n   t h e   F i l e   C h o o s e r   c h a n g e s   t o   t h e   s e l e c t e d   d i r e c t o r y .   
--IJHG @ �  Ld
   �kt P  LNOMLQTRT!	  M a r k P r o c
C  � U n m a r k P r o c
a  � H i s t o r y M e n u
�   � WXVU` | X !	ab`_ \][Z"&  ��	((e"a { H i s t o r y   M e n u 
 
 U s e   t h e   H i s t o r y   M e n u   t o   q u i c k l y   n a v i g a t e   y o u r   f i l e   s y s t e m . 
 
 T h e   H i s t o r y   M e n u   c o n t a i n s   t h e   f o l l o w i n g   t w o   s e c t i o n s :   H i s t o r y   L i s t   a n d   M a r k e d   D i r e c t o r i e s   L i s t . 
 
 H i s t o r y   L i s t 
 
 T h e   H i s t o r y   L i s t   l i s t s   t h e   m o s t   r e c e n t l y   v i s i t e d   d i r e c t o r i e s ;   u p   t o   f i v e   d i r e c t o r i e s   c a n   b e   d i s p l a y e d . 
 
 I f   y o u   v i s i t   m o r e   t h a n   f i v e   d i r e c t o r i e s ,   t h e   o l d e s t   d i r e c t o r y   i s   r e m o v e d   f r o m   t h e   b o t t o m   o f   t h e   t h e   l i s t   a n d   t h e   n e w e s t   d i r e c t o r y   i s   i n s e r t e d   a t   t h e   t o p . 
 
 T h e   H i s t o r y   L i s t   i s   s a v e d   f r o m   o n e   e d i t i n g   s e s s i o n   t o   t h e   n e x t . 
 
 M a r k e d   D i r e c t o r i e s   L i s t 
 
 T h e   M a r k e d   D i r e c t o r i e s   L i s t   c o n t a i n s   d i r e c t o r i e s   t h a t   h a v e   b e e n   m a r k e d   f r o m   t h e   S p e c i a l   M e n u .   M a r k e d   d i r e c t o r i e s   p r o v i d e   q u i c k   a c c e s s   t o   f r e q u e n t l y   u s e d   d i r e c t o r i e s . 
 
 M a r k e d   d i r e c t o r i e s   r e m a i n   i n   t h e   H i s t o r y   M e n u   u n t i l   y o u   u n m a r k   t h e m .   T h e y   a r e   a v a i l a b l e   f r o m   o n e   e d i t i n g   s e s s i o n   t o   t h e   n e x t . 
 
m T o   u n m a r k   a   d i r e c t o r y : 
 
 1 .   N a v i g a t e   t o   t h e   m a r k e d   d i r e c t o r y . 
 
 2 .   S e l e c t   U n m a r k   f r o m   t h e   S p e c i a l   M e n u . 
 
 T h e   d i r e c t o r y   i s   r e m o v e d   f r o m   t h e   M a r k e d   D i r e c t o r y   L i s t   i n   t h e   H i s t o r y   M e n u .   
 d $  "� S p e c i a l   M e n u 
 
 U s e   t h e   S p e c i a l   M e n u   t o   d i s p l a y   y o u r   h o m e   d i r e c t o r y   o r   t o   M a r k   a n d   U n m a r k   d i r e c t o r i e s . 
 
 T h e   S p e c i a l   M e n u   c o n t a i n s   t h e   f o l l o w i n g   t h r e e   i t e m s :   H o m e ,   M a r k ,   a n d   U n m a r k . 
 
 H o m e 
 
 S e l e c t   t h i s   o p t i o n   t o   d i s p l a y   y o u r   H o m e   d i r e c t o r y   i n   t h e   F i l e   C h o o s e r . 
 
 T h e   H o m e   d i r e c t o r y   i s   a   d i r e c t o r y   d e s i g n a t e d   o n   y o u r   s y s t e m   a s   y o u r   s t a r t i n g   p o i n t   f o r   f i l e   o p e r a t i o n s . 
 
 M a r k   a n d   U n m a r k 
 
 U s e   t h e   M a r k   a n d   U n m a r k   o p t i o n s   t o   a d d   o r   r e m o v e   d i r e c t o r i e s   f r o m   t h e   M a r k e d   D i r e c t o r y   L i s t   i n   t h e   H i s t o r y   M e n u . 
 
 M a r k e d   d i r e c t o r i e s   a r e   d i r e c t o r i e s   t h a t   y o u   m a y   w a n t   t o   a c c e s s   q u i c k l y   o r   f r e q u e n t l y . 
 
� T o   m a r k   a   d i r e c t o r y : 
 
 1 .   N a v i g a t e   t o   t h e   d i r e c t o r y   y o u   w a n t   t o   m a r k .   
 
 2 .   S e l e c t   M a r k   f r o m   t h e   S p e c i a l   M e n u . 
 
 T h e   d i r e c t o r y   i s   n o w   m a r k e d ,   a n d   a p p e a r s   i n   t h e   M a r k e d   D i r e c t o r y   L i s t   i n   t h e   H i s t o r y   M e n u .   
� V i e w   M e n u 
 
 U s e   t h e   V i e w   M e n u   t o   s p e c i f y   t h e   o r d e r   i n   w h i c h   t h e   c o n t e n t s   o f   a   d i r e c t o r y   a r e   l i s t e d   i n   t h e   F i l e   L i s t . 
 
 T h e   c o n t e n t s   o f   a   d i r e c t o r y   c a n   b e   s o r t e d   b y : 
 
 * 	 N a m e 
 
 * 	 D a t e   M o d i f i e d 
 
 * 	 D a t e   C r e a t e d 
 
 
 j  fged%> "lkljio (  = F i l t e r s   M e n u 
 
 U s e   t h e   F i l t e r s   M e n u   t o   s p e c i f y   t h e   t y p e   o f   f i l e s   t o   l i s t   i n   t h e   F i l e   C h o o s e r . 
 
 T h e   F i l t e r s   M e n u   i s   n o t   a l w a y s   a v a i l a b l e   i n   t h e   F i l e   C h o o s e r . 
 
- V o l u m e s   M e n u 
 
 U s e   t h e   V o l u m e s   M e n u   t o   s p e c i f y   a   d i s k   l o c a t i o n   t o   s e a r c h   f o r   f i l e s . 
 
 T h e   V o l u m e s   M e n u   i s   n o t   a l w a y s   a v a i l a b l e   i n   t h e   F i l e   C h o o s e r . 
 
 
 
n  t  pqon)� "yuvts= A r r o w   B u t t o n s 
 
 U s e   t h e   A r r o w   B u t t o n s   ( t o   t h e   l e f t   o f   t h e   F i l e   L i s t )   t o   m o v e   t o   t h e   d i r e c t o r y   i m m e d i a t e l y   a b o v e   o r   b e l o w   t h e   c u r r e n t l y   s p e c i f i e d   d i r e c t o r y . 
 
 
y &� x "z{yx � P a t h   P o p - u p   M e n u 
 
 T h e   P a t h   P o p - u p   M e n u   i s   l o c a t e d   a b o v e   t h e   F i l e   L i s t .   T h i s   m e n u   d i s p l a y s   e a c h   d i r e c t o r y   i n   t h e   c u r r e n t   p a t h . 
 
 T o   d i s p l a y   t h e   c o n t e n t s   o f   a n y   d i r e c t o r y   i n   t h e   c u r r e n t   p a t h ,   s e l e c t   t h e   d i r e c t o r y   f r o m   t h e   P a t h   P o p - u p   M e n u . 
 
 F i l e   L i s t 
 
 T h e   F i l e   L i s t   l i s t s   t h e   c o n t e n t s   o f   t h e   c u r r e n t l y   s p e c i f i e d   d i r e c t o r y .   T h e   i c o n   d i s p l a y e d   b e f o r e   e a c h   n a m e   i n   t h e   l i s t   i n d i c a t e s   w h e t h e r   t h e   l i s t i n g   i s   a   f i l e   o r   d i r e c t o r y . 
 
 U s e   t h e   F i l e   L i s t   t o   s p e c i f y   a   d i r e c t o r y   o r   f i l e   f o r   t h e   c u r r e n t   o p e r a t i o n . 
 
 
} ,  � P a t h   N a m e   T e x t   F i e l d 
 
 T h e   P a t h   N a m e   T e x t   F i e l d   d i s p l a y s   t h e   n a m e   o f   t h e   f i l e   o r   d i r e c t o r y   s e l e c t e d   i n   t h e   F i l e   L i s t . 
 
 U s e   t h i s   e d i t a b l e   t e x t   f i e l d   t o   s p e c i f y   t h e   p a t h   n a m e   o f   a   f i l e   o r   d i r e c t o r y . 
 
 
 
~  �� �~} � C o n f i r m a t i o n   B u t t o n s 
 
 U s e   t h e   C o n f i r m a t i o n   B u t t o n s   t o   a p p l y   y o u r   s e l e c t i o n   i n   t h e   F i l e   C h o o s e r . 
 
 
 
-� ������ ��"a�  ��  ���� �0   5j/�8  P a t h M e n u
.�    F i l e L i s t
.� 	   � -
	
 &(,.                                             i R e s i z i n g   t h e   F i l e   C h o o s e r 
 
 M a k e   t h e   F i l e   C h o o s e r   w i d e r   t o   d i s p l a y   u p   t o   f i v e   d i r e c t o r y   l e v e l s   a t   a   t i m e .   T h e   c u r r e n t   d i r e c t o r y   i s   a l w a y s   d i s p l a y e d   i n   t h e   l e f t m o s t   l i s t .   A d d i t i o n a l   d i r e c t o r i e s   c a n   b e   d i s p l a y e d   a s   f o l l o w s : 
 
 * 	 C h a n g e   t h e   c u r r e n t   d i r e c t o r y   w i t h   t h e   P a t h   P o p - u p   M e n u .   T h e   n e w   c u r r e n t   d i r e c t o r y   i s   d i s p l a y e d   i n   t h e   l e f t m o s t   l i s t   a n d   t h e   o t h e r   d i r e c t o r i e s   i n   t h e   p a t h   a r e   d i s p l a y e d   i n   t h e   r e m a i n i n g   l i s t s .   T h e   d i r e c t o r y   n a m e s   a r e   d i s p l a y e d   i n   t h e   t e x t   f i e l d s   a b o v e   t h e   l i s t s . 
 
 * 	 S e l e c t   a   d i r e c t o r y   f r o m   t h e   F i l e   L i s t .   T h e   c o n t e n t s   o f   t h e   s e l e c t e d   d i r e c t o r y   a r e   d i s p l a y e d   i n   t h e   l i s t   i m m e d i a t e l y   t o   t h e   r i g h t ;   t h e   s e l e c t e d   d i r e c t o r y ' s   n a m e   a p p e a r s   i n   t h e   t e x t   f i e l d   a b o v e   t h e   l i s t . 
 � 	AttributeContextqBlock!untQsExtraKeywordBlockLengthasinkListAType	NodeBlockADataA	TextsOffsetasTagextAAttributes	itleQs
ypeVersionvhelpDocument<�    |  �    j r0m�k                                                                                                                                                                                                                                                                                                                                                                         q 2 �qb b!qb6b �B
yarVAb/!qNbaaI"Eqb,(qbK&q."�&!;bo&qEb�&!Kr,&qSb�&aYr�&a^b�&acr#�&qh"#�&qmb&�&!rb&�&aw"'�&a|b-�&R �.�"& �r.�&ar?aq!buq!%bGbTr,"�r,"�r,"�b,"b,"=b,"[b,"yb,"�","�b,"�b,""(3b,"�r""cb+b.<b,4h",4�b,4�2,4�,4;b,4[r(wb,4�bfbb�r_r;�b,A�b,A�R,A�rn,aAr�Qbcab�ar�ab�(abarq"!b�qbaKb4,aP"V,aP"�ar,qPrxar(ab�qb>ar:q"�qb�ar�q"�!r�!r�a"�a"�qr�qb�ab�ab�ab�ab�!b�qr#�Qb#�ab#�ar#�q"#�ab#�ar#�ab&qab#�a"&l!r&�!r&uq"&�ab&�!b&yqb'�ab&}ar'�!'�R'�ab+�a"'�qb-�ar+�ar-�!r.z!B-�a".�qr.�Qb-�(ab.�ab.�!b.�qb.�qb.�b �.�b, �b.��   r, �r/�