��     	  �d  � S e t C o l o r  S t y l e   C h o o s e r"kg   $ T h e   S t y l e   C h o o s e r�'>�� ��  ��   ��   ��   ��   ��   ��   ��   �� 	  ����& S t y l e   D i s p l a y   A r e a$ A t t r i b u t e   T o g g l e s& S p e c i f y i n g   a   S t y l e X � �Sbs��� A s c e n t D e s c e n t F o n t   S i z e  S e t   F o n t   B u t t o n" S e t   C o l o r   B u t t o n* C o n f i r m a t i o n   B u t t o n s O v e r v i e w�# A^u����� S i z e F i e l d"`8I S p e c i f y S t y l e s A t t r i b u t e s" S t y l e D i s p l a y A r e a C o n f i r m B u t t o n s A s c e n t F i e l d S e t F o n t v s t y l e c h s r D e s c e n t F i e l d    *  �� s t y l e   c h o o s e rJ<"%+09?DINS   & !"#$ S p e c i f y S t y l e s' 
    (" S t y l e D i s p l a y A r e a
�    � A t t r i b u t e s
�    �+ S t y l e   C h o o s e r 
 
 U s e   t h e   S t y l e   C h o o s e r   t o   s p e c i f y   s t y l e s   f o r   s e l e c t e d   t e x t   i n   a   t e x t   f i e l d . 
 
 T h e   S t y l e   C h o o s e r   c o n t a i n s   t h e   f o l l o w i n g   c o m p o n e n t s : 
 
 S t y l e   D i s p l a y   A r e a 
 A t t r i b u t e   T o g g l e s 
 S e t   F o n t   B u t t o n 
 S e t   C o l o r   B u t t o n 
 A s c e n t   F i e l d 
 D e s c e n t   F i e l d 
 S i z e   F i e l d 
 C o n f i r m a t i o n   B u t t o n s 
 
 
 S e t F o n t
,    � S e t C o l o r
H    � A s c e n t F i e l d
f    � D e s c e n t F i e l d
�    � S i z e F i e l d
� 
   � C o n f i r m B u t t o n s
�    �(  5   )*('  ))(��   O O O � � � �-��./-,"aV!       6:78  ��!V
  LL3421  
�   �; A t t r i b u t e s
�    �< "� A s c e n t F i e l d
	6   �
	Q   � 5 S t y l e   D i s p l a y   A r e a 
 
 T h e   S t y l e   D i s p l a y   A r e a   d i s p l a y s   a n   e x a m p l e   o f   t h e   c u r r e n t   s e l e c t i o n .   A s   y o u   c h a n g e   y o u r   s e l e c t i o n ,   t h e   c h a n g e s   a r e   r e f l e c t e d   h e r e . 
 
 
 D e s c e n t F i e l d S i z e F i e l d^  B  =><;  "BCA@� F o n t   S i z e 
 
 S i z e   r e p r e s e n t s   t h e   s i z e   ( p o i n t   s i z e )   o f   t h e   f o n t . 
 
 T h e   f o n t   s i z e   i s   i n i t i a l l y   s e t   t o   " A u t o " - - t h e   d e f a u l t   v a l u e   s p e c i f i e d   b y   t h e   a p p l i c a t i o n . 
 
 T o   r e t u r n   t o   t h e   d e f a u l t ,   c l e a r   t h e   f i e l d   a n d   r e a p p l y   t h e   s t y l e . 
 
 
E 	� F "	 L  GHFE� "LMKJO    P  VTQRPO VWUT b!��$                        ] A t t r i b u t e   T o g g l e s 
 
 U s e   t h e   A t t r i b u t e   t o g g l e s   t o   s p e c i f y   t h e   f o l l o w i n g   s t y l e s : 
 
 B o l d 
 I t a l i c 
 U n d e r l i n e 
 H i d d e n 
 S t r i k e t h r u   
 
 T h e s e   s t y l e s   a r e   s p e c i f i e d   w i t h   t r i - s t a t e   t o g g l e s .   T r i - s t a t e   t o g g l e s   h a v e   t h r e e   s t a t e s :   
 
 S e l e c t 
 T h e   s p e c i f i e d   a t t r i b u t e   i s   a p p l i e d . 
 
 U n s e l e c t 
 T h e   s p e c i f i e d   a t t r i b u t e   i s   r e m o v e d . 
 
 N o   S e l e c t i o n   ( " F u z z y "   S t a t e ) 
 T h e   s p e c i f i e d   a t t r i b u t e   i s   u n c h a n g e d   w h e n   t h e   s t y l e   i s   a p p l i e d . 
 
 
 S e l e c t i n g   t h e   F o n t   a n d   C o l o r   t o g g l e s   e n a b l e s   t h e   S e t   F o n t   a n d   S e t   C o l o r   b u t t o n s .   S e l e c t   e i t h e r   o f   t h e s e   b u t t o n s   t o   o p e n   a   c h o o s e r   t o   s p e c i f y   f o n t s   o r   c o l o r s . 
 
 
 
� A s c e n t 
 
 A s c e n t   i s   t h e   s p a c e   a b o v e   t h e   b a s e   l i n e .   S p e c i f y   a   v a l u e   f o r   a s c e n t   i n   t h e   A s c e n t   f i e l d . 
 
 A   l a r g e   a s c e n t   v a l u e   i n c r e a s e s   t h e   d i s t a n c e   f r o m   a   l i n e   o f   t y p e   t o   t h e   l i n e   a b o v e   i t . 
 
 A s c e n t   i s   i n i t i a l l y   s e t   t o   " A u t o " - - t h e   d e f a u l t   v a l u e s   o f   t h e   f o n t   a r e   u s e d   f o r   t h e   a s c e n t   v a l u e . 
 
 T o   r e t u r n   t o   t h e   d e f a u l t ,   c l e a r   t h e   f i e l d   a n d   a p p l y   t h e   s t y l e . 
 
 � C o n f i r m a t i o n   B u t t o n s 
 
 U s e   t h e   c o n f i r m a t i o n   b u t t o n s   t o   a p p l y   y o u r   s e l e c t i o n . 
$`   ^pb� ``!aaQ(Qawz2b2D&                                     � T o   s p e c i f y   a   s t y l e : 
 
 1 .   I n   y o u r   a p p l i c a t i o n ,   s e l e c t   t h e   t e x t   y o u   w a n t   t o   s t y l e   o r   p l a c e   t h e   i n s e r t i o n   p o i n t   w h e r e   y o u   w a n t   t h e   n e w   s t y l e   t o   b e g i n . 
 
 
 2 .   F r o m   t h e   S t y l e   C h o o s e r ,   d o   a n y   o f   t h e   f o l l o w i n g   t o   s p e c i f y   a   s t y l e : 
 
 * 	 S e l e c t   ( o r   u n s e l e c t )   a n   a t t r i b u t e   t o g g l e . 
 
 * 	 S e l e c t   t h e   F o n t   t o g g l e   t o   e n a b l e   t h e   S e t   F o n t   b u t t o n .   S e l e c t   t h i s   b u t t o n   t o   o p e n   a   F o n t   C h o o s e r . 
 
 * 	 S e l e c t   t h e   C o l o r   t o g g l e   t o   e n a b l e   t h e   S e t   C o l o r   b u t t o n .   S e l e c t   t h i s   b u t t o n   t o   o p e n   a   C o l o r   C h o o s e r . 
 
 * 	 S p e c i f y   t h e   A s c e n t ,   D e s c e n t ,   o r   S i z e   f o r   s e l e c t e d   t e x t   i n   t h e   a p p r o p r i a t e   f i e l d s . 
 
 T h e   S t y l e   D i s p l a y   A r e a   d i s p l a y s   a n   e x a m p l e   o f   t h e   s p e c i f i e d   s t y l e . 
 
 
 3 .   A p p l y   y o u r   s t y l e   w i t h   t h e   c o n f i r m a t i o n   b u t t o n s . 
 
 T h e   s e l e c t e d   t e x t   c h a n g e s   a c c o r d i n g   t o   y o u r   s t y l e   s e l e c t i o n s . 
 
 
 
� S e t   F o n t   B u t t o n 
 
 T h e   S e t   F o n t   b u t t o n   i s   e n a b l e d   w h e n   t h e   F o n t   a t t r i b u t e   t o g g l e   i s   s e l e c t e d . 
 
 S e l e c t   t h e   S e t   F o n t   b u t t o n   t o   o p e n   a   F o n t   C h o o s e r .   F r o m   t h e   F o n t   C h o o s e r ,   y o u   c a n   s p e c i f y   a   t y p e f a c e   a n d   f o n t   f o r   y o u r   s t y l e . 
 
 
u                                                                                                                    � D e s c e n t 
 
 D e s c e n t   i s   t h e   s p a c e   b e l o w   t h e   b a s e   l i n e .   S p e c i f y   a   v a l u e   f o r   d e s c e n t   i n   t h e   D e s c e n t   f i e l d . 
 
 A   l a r g e   d e s c e n t   v a l u e   i n c r e a s e s   t h e   d i s t a n c e   f r o m   a   l i n e   o f   t y p e   t o   t h e   l i n e   b e l o w   i t . 
 
 D e s c e n t   i s   i n i t i a l l y   s e t   t o   " A u t o " - - t h e   d e f a u l t   v a l u e s   o f   t h e   f o n t   a r e   u s e d   f o r   t h e   d e s c e n t   v a l u e . 
 
 T o   r e t u r n   t o   t h e   d e f a u l t ,   c l e a r   t h e   f i e l d   a n d   a p p l y   t h e   s t y l e . 
 
 
 
 � a-q!!
aqaa!!a	
aaaaaq!Qaqaq!aqaa!
! &
qa!(aqqa,q!x                                                                                                                       � S e t   C o l o r   B u t t o n 
 
 T h e   S e t   C o l o r   b u t t o n   i s   e n a b l e d   w h e n   t h e   C o l o r   a t t r i b u t e   t o g g l e   i s   s e l e c t e d . 
 
 S e l e c t   t h e   S e t   C o l o r   b u t t o n   t o   o p e n   a   C o l o r   C h o o s e r .   F r o m   t h e   C o l o r   C h o o s e r ,   y o u   c a n   s p e c i f y   a   c o l o r   f o r   y o u r   s t y l e . 
 
 
 � aqa!	AttributeContextaqBlock!untaQsExtraqKeywordBlockqLengthaasinkListaATypeq	NodeBlockADataA	TextsaOffsetqasTag!extAAttributes	itleQsa
ypeVersionavhelpDocument`                                                                                                                                                                                                                                                                                                                                                              � 1W@bDr<b �b
Gq"8ar
qr"a!Lb �b �bQb(jr&%B&+F"&0�r&9	zr&?	�b&Dyb&I�"&N�b&S�b&^R}q"Ma"Iq"fars,qr�,a"�,!b=,a"[,Ab,!B�,ar�,!"�aaP",�"�r�b�r�bb-rbN"Wb(blbzbsb�b0er,5�b,5�,�5�b	fb,5�"r��"�"	�b	mr	�b	�"	qb\"	ubhbWbcb�blb�b�"pr�bt"�b�r�b�r�b�b�b�B